# ====================================================================
#
#      altera_avalon_cf.cdl
#
#      Configuration file for the Altera Avalon Compact flash driver.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####

cdl_package CYGPKG_ALTERA_AVALON_CF {
    display       "Altera Avalon Compact Flash"

    parent        CYGPKG_IO_DISK_DEVICES
    active_if     {!CYGHWR_DETECTED_SOPC_DEVICES || is_substr (CYGHWR_DETECTED_SOPC_DEVICE_LIST, " altera_avalon_cf ")}
    active_if     CYGPKG_IO_DISK

    description   "
           This option enables the compact flash driver."

    compile       altera_avalon_cf.c 
    compile -library=libextras.a altera_avalon_cf_devices.c

    cdl_option CYGPKG_ALTERA_AVALON_CF_CFLAGS_ADD {
        display       "Additional compiler flags"
        flavor        data
        no_define
        default_value { "-I`cygpath -u $$SOPC_KIT_NIOS2`/components/altera_avalon_cf/inc -I$(PREFIX)/include/cyg/hal" }
        description   "
            This option modifies the set of compiler flags for
            building the Altera Avalon compact flash driver.
            These flags are used in addition
            to the set of global flags."
    }

    cdl_option CYGPKG_ALTERA_AVALON_CF_CFLAGS_REMOVE {
        display       "Suppressed compiler flags"
        flavor        data
        no_define
        default_value { "" }
        description   "
            This option modifies the set of compiler flags for
            building the Altera Avalon compact flash driver. These flags are removed from
            the set of global flags if present."
    }

    cdl_option CYGDAT_ALTERA_AVALON_CF_SECTOR_SIZE {
        display       "Disk sector size"
        flavor        data
        default_value 512
        description "
        This option controls the disk sector size (default=512)"
     }

    cdl_option CYGDAT_ALTERA_AVALON_CF_USE_MBR {
        display       "Use Master Boot Record"
        flavor        bool
        default_value 1
        description "
        Expect the first sector on the device to contain a master boot record."
     }
}
