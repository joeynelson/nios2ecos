��/  �d>$Lw�e�,]�b�sᗸ@[����h/m<�=O�����M�XX�+�*�Ͷ�����,��8K���y݋N��T��c�����aQ�h/����M{����Qe$�q�Hw�.�6n���@bJK;˵�泿�
��=$=�K�V�&��6`�St�fd��B�Ã֧��O"�CR��c(^�!�~W����B����Y��g��A�y[3Ղ�㲕�������ч�/tsn3������G"�bb��fu2%P ��ڹh:�~9CG��ߤ������H,��!әj�q�
5-����g`Hv���Q�<�ZR��v�����C@kl��~1>"i��b�aް��X��9U���-�ÿ�GO/1��*��04j�vQDU�J�����B�₨>��q�5,�O>��L�֡�<��P<Å 2<uwY����Ğ�O�C���-Li��bRԡ�r���ƨ�"��4�V*m[���D�+�K����4��MB�@Q�J}��P��5�tG����h�ݟv�/&�(d=�+o_@ ���U��$M��2��:E��պ2�꯷p��\�sD�bWY����	*��s��9��u�,�L��w��N���j�~�v�N׺�,E�V�[cCR&>k���dh��WQx����ǎ	���`xW�
���g��g�}�|%�f���ҙ[�C�a*kk�ѳ�n����	�
�9�J�
[>e���ӎ��*���t��ʶ������ΉsloBJn�K�tr(~ܯq�DOV3Ϳ�qߢ�k��@�H%"�
�$��U?��^�\k��eֹ:����0n�=}������f�I7?0�g^�֎j�a�⟍�N�����I!?ɰf���e`:��Ew�UԡO�\�#��!q?j���hoaf���������)ۃ��>Dt-�z��a�2�%����Mh��a���3��]�����g�䌓ɨ#K��خ*�a�'���	�����i�����]sq�p�<kH=d��V eJ�D��r�(��bm��?�/���3��>��AB�k����S7|�����G�"iw�eФC���$��Jd�`�~�U��&;" �W[�~�ru�Pa@Y��9�ǈ^�w�����=��p:�IjᏅ����[1x�a�:,�}]��3�o�%!��z f��Y�B�U��?�l�Q�I��J4�e�BH��x��o6u���8��`��7n	���X��A%6�=���I ����A�k�!$��}=fFC0$z�w%J1ےLn�L-�[��%�_vwޕ�|�^̸� ����?�y��O���<���qU_D����P��Z,>]����E}��,��+��Б�n�ڍ^��8c_������f@}`-C����.')���֖�5�!B���p�*��������6�X: V�%h���2?Fr��`Hr��8�Ez;Λ�\��"x�k�K�?�Q�N���k&ބ�<�K�0G��O��Q�v�O�ؼ�y�8��'��w�J@P��8I��FK���?���Dl7���޼f�ϖ�s5bK͆D{�"��>�*��v��$1z;�6?z4��}�y�B�\:tE�2�k�{��o>e~�š�
�O�G��[�h�<&��:�=��m�}],%dmjj��B�Db֫F�:�]qo��68�����$��N����/&��fɋ#�?��?��r����k�m�D�VhOoߋoĶ��a/�s����,=��yZ�Ӹi�[��\C��G�c�.�ѧ7_�DOJ}(��ux���Ҿ�(�-��o��SAUe�e���1a��88o�/�=خ�u2�P��u~�,�[Q5��C��U�5Y��N�0=���Ϭ'���yY! Q��)�$�}��#��:	u�TN��\݈9�=�n'�����N1^z�D
J�eiv�7��d�������[-�hfD.�32l鸵�)fys#�9Q~����ͽ	���R��`���bĩ�㷲�򕗪�F![2�8�Y`�|�n8z�Y&�ҷ�yl�Laj����̔� ?��.ҐLk���y6�wE���f],�����B�`z�.�p|��|���,W�4xt�$�#YO�CIGhz�b0���(u�ɸȵ= ��?�2M8�Z#�ϰU�!�)�mmn�J�$�΄�淢�L�7G4�vP�gt������O,�a�;v;��]R��;-��PSAe$uU��Nr���~�&�xR�$���ͺ��E}1�/�ȉ��S����D ���xS&a�/�q�{��?�v����y���������"l4���*���6h�-y����(�i��~g�])��o��`��)8FEJ�D�l*�ǀV�l�A���{�AF�ra�&�"���,ޠ��X!��O�Y�P%@�RVA�=� Z�g��?)�#�9$@``t3'�	s����9��F��ޖO�+�a��� T5�%����dG,��1!ѣ� � :��	�X`�,O��F�?�g��TR)����$�!{���5��TF����;?9�}�hڱտ��9����#o&dQ��) ��V�x~M3�mb���������'��^V�	)�v唛���%�s!�v�JYA����G9S��`�^��q��Z�TǮ o��9�[���<+�����<���|[	X(K+��CJTvML4AW�(t:�:�B}?ǥw�����y~�DXP��\(�:r뜭Y裬c�ND&��Ĩ��B��n�Ek(�,��:�}m�雙�*I�V:#���Q�=c��Cɇ!S(���J���\%�''����__�%4�!������B7�չ�7�\C���CCIF$���1s�-.��@�K��j��$�r�4��r�����|1���1{��M戻��<�w7f���gV.0�z!���J�RJ#��5X��u�`�,������W^�co�
�gZ'i�>ճ르�:��'�I��)O�d�ԏ1m��,ƚ���7M7��{JJ/L���j��թkR�,�[���� �E�ڱ/������kIdoJ�.S�����3���y�Q�6��2?=Mi���<V�Dx�����}0����@B]`Nѭge��y	�	��$hRJ�X(aT�G]j�#���4gu�U���Ҙ�s~A.�]�T�|�)�ي�X�ʄ�Qމ��9��0�e�D�^U:�Xg�����n��B�u'�N^�M`�؂�D¨ҿ����Nx��=G%��~�l�����a:��o�T���=�7-��4�m�`8�ڥ�u��14}�DXK�':��u�I�Sڐ7���f��+U���k���e�3����11�fV���	�SY�Qw��;,TH\c��HNBZ�?����?E!�z�͹R�U�k�k}�3KDf"��z"U���d����,��Gc.���EG���~���`bQ��<��|(�G�1�$˨��NU���V.0�dg��C=��S3�	��B��;�ZH���྄�)[��A=/��]ZM�lt�C��:R2�n�/	��<�f�D�Q'�afa߰�ה�m��df�[1�W��F���jx���ʟ#"|�;�i�6���){��9�~� ���;�����Hh6g��f9wI1�.�i<w�'�,#Q��Lo��5>
��4r�z?(C�uyk�p��(��Z�WY�7�����޿�g�_����6*����6 ���Y�ޔetߺ����׀K/v*���4��ߺ����y���H�q(rJ�:]���קYߒ'����"W���٨��d�|��܅7V���R����DA��_�m���/�V�5�rV�ռ�7�y��v��It����Cַ`�ȧs�VV3|9d��I�˜	���y�)FoHb��f�d��/P�0���M�g�*�@��,�����K�}���}��
o������}&v�Ł2$'̉��Y9�M�u�x�x.�C�}c@d$�L�RF�23)�=L��B�o��^�H�;�4[�ɂ�s�L�f	s�0�@xZ���8�J�>�y�K�����.��;����5���a��%���5�b�6�}�Co|��q�w��]�ߏfi3�����17+�l�K.�R�I���g�=�V)�d�O0C04�&��δU?7EC�O9m����G�F��E\~���m�.�6XP�Y�[i��6A-�t�,M������紎��j�8�w)iB��M^Z���K��C�gۊF&G��j�+�ʛ���(y�4'�N�Y�w��CRs��-R�S���~l���CR�kO��8f�_���t���I �4�*݄�-����J�+��kXn�S��8	w��w�v3���H�W� 2�S�Fk�^���;!�Y����Z��#��9B8����bE���2L艛���q���%R:a�kiq���J���$�`{Fh��u-�5��+���%4����=�\�P����,��bM	��cւY�GVyCL3�C!�����1��њ�!��UV��#�P�����xQ�HKV�{I�gd�1�o�{�T�v��ps�2
�5���������y��b�+^3�
2����ت[#������x��CJ���3�"�QRa��d��^SД���U�tȧB�b��э���IN#����oswډE�c��+��r����|%|�,�J�� �2�ın��=� ���H琢=Ǹ-�U	s"4غO}�G��O���嵃fj�ݝæ�^$�Q>lԎ�y$6�}2e����hj \s[�E]$�h �h�K���ȼKL�[1���v7|sۨeى�b����kӑ��������f����z��Ѽ~�EWZ�����Ň
�ax�;^��妴��O���܆����7�b2sPt	��r�rjV�Rؕգ.D_���h�|7a�X9�G�ܰ+��{Fވf���)l�]F��f'�biM���5�_�/�,���I����S�������&劻*B�<�	�J��J�d;�%�uę5#��%pl9��ݶ\���P����.hl�.,v
P�ꓽ�M�6�+K��p�"�8�o��ݙ��C�X5�i@i�4�,~���	276���l��_:U��[��B��WW1Y����&�)�:�o�쳸��ʢKx��˶W�U���z�E�����lF�,�^g4�v���?O��̞f�[wWJV&�N(��X�������%��y��_���@�����$��ݒB��ѫd�an�;q��r^�a�.?*'sJ�Q��=��s�_um���� ,�mq�6^���k\�8�%����YF[q�Z1b�X1���S"��yPoZ|y;��J�l����w.�r���:�#ir��8|����/TЀ,�ʆχ�	y}B��&��v7͗�&Dc�bu���_ud��K�c!��c�O�I�LG�����r�)�z�TsЉ�Y�?��P��	��3yt�Ͼ��+D�v�M��h��kx�o�� 0'��MЛ���"�T�٘�Ŗq��ɔ$��y�2b�bk�x;ʨ(ƤH��,K�ܠ�0D�ت.K�����,��߀�5b����(溮����JZS�F]h�������f�������3��gǪF/��-�������c�05�UFs#K��L�C���C�<�b9�墈y�t�R����u��X�)	ڳQ�j^YQ��1�ln�����S;"e���/�Ñ�ExBe�����ύj��O��S>?y(�'�EU(vz�c��ڇ#�ef�@Z�e[
 �e�?��W�=W�?�AЬ��S@)��"��rՠJ�wk��3C��-3	L�&���t_;��u�t`����B��;�f��g�k���ƥF�l�1��}|@��怐�pokȺl�����"��yGw�I�6"k�5��f�KYg7��-/$��c0�<;�*�i�6�9����4E�W�k�wSS����b��V�Lc�l���=��]�b���;0n�)4�O�u�a��d�v�fVt� ����S�H�i����a�8���P���YD:��²-B������6W�Iu7|`��-Me�eu���9���l�z�5^��h��f�
з�=L�g�D�)�l��\e�歃��J.d�O�wC��e>�E#�wS���|�<dEf�u[8|��2�d<EBT*R6j�
V�*6�Z�M`k��B�z�*:�V!	�$F�v�A\R�t��,��Y��z�Ad��FEу�!Ɓ�׶���4��w��
�ly����~�.���vȑ@�9�#|M�y|Ra�"HN������8�V��X�9���^n�I�E�x�3�i�x[�MK��=a�0�}�5�1x������Xů�.�@���?�@{c���x�R�9��8�-|��jr��`1��h���QIE�����Y'xտꔵ������[��"����CT�k��A��{;9�SU�af��4�,K?n�b�T_��4i�b1s�t�·���@�����-_/��"�����7܃F�#�YZ��߰2��h8܎��So���3&Ek0��~�Ͻ�H�-ƱglW��ɋr!��A�`rЬ���Z4O��f����w�;�	�q�/����H�<o�ƃ���R�nsβӢ�`�s����ZO��K� C]k�*B=�Q�=�m��R��g�t����z	�'���� ��\f�3�����=nY&���DLO���Y:��d�"���)�����2�;�؃5Z�REG�&ig�4�1�≵�����H�J� ^������SwW�����T�H$����9�T�U��
t�N-w�2v�ffM��v�0�v��ޒ�t��o��e��;HWs�-\��(����_�`����+7Z��Ԙw��K�X{%{���JuUʬ��9�����"���W��R��R�&pc�K[��\�ʏo�sn�d�Z��4"Y���+�ɞ����C")0��gO푸��G�i���3L��	Y�7�>������Ué�K�%�QR��z.�1��X(�KU�!���,j.�������;�tѬ'���x9Hw&V��?��_��!��W��w�a�(>��'�+�x�³2���0JN36������IC�!�.�n>��$Q@���~�LI�A��R�Kb�޲!����N/W^����㏀�*.����ui�s���;hvlh���Ǉ�i%���:��)���l�p�����[����GW�֩��Ϣ�a��9BbKk0�&ZE8�������Wq^�Y�"��1��R�,�gu�V�寈B0A/p�s����*�鏟����}����lA�y?������y�~}�h�3^�@,:h��0޿Y�$p�R�����N��i�2�= ��?�~^v����d&ȝ7���^g��Ky��� t���Yp�G�!�7Ҵ�&�V}�	aԤ�B}� E�4~Z�H6NX7�/]�팞<�1yT4�Q��Y�Cn�O�߱ѺD,M�&���X|�@*�뷝Ԩ����g����FįZOa���V�2I33;����(�u�ɰ��ƴ�f�/zdw��R�dOnj�2+.��/�O؇Wsk1#LR�he ��b+��M�_��	|�t1�ky�D���+����&&U��  �f.��R�lDK, Q����%@	D��j�v���Y�"E��_�Ğ�
�I"n�Rx�:#%S�[�����pi�C��i���ŦN\�/;��s��NYj>h|��ԐEtT���ԩt�����Z����_�`V�;'��gI`Y�L��=�Nl'a�h)cc�R�W�s$���.���!�$���R8� _H�HR-O~��?�T�5��2Ep�פ���C+*2x��"�x�/�=���t�"L!����ǲ�"ϕ��@p$9�D<��D,_ǉ�y�5�������6��2���P�F2�p����n�xF�B덀��n�gZwfգ��"Gj<� �88�{�e����O<|$�H�G�Om:p���@#q�ܢ\4�"� &�ߺ�D�,o��?y!�9#a��7�Y���T�����0�X�6��D\)����T�� e�����ĉh_4�Ѩ�va��~�X�h�N`ޖte!��.|�bX�ˈ��|��,������ -�Srt���J�� ��~� �̝#�����w�чR�C^�֔��=�#s��ut6Hmk���,(j�@�桯cxN���p�������HP��Mt�Y,�Al=v�c��yǱ�y�e?�aW0;�14,b�Y�x�NI���K.$�kd��̫��S�n%\A9j7��6#�Z�=���!��v�>	:�<�l�oލ2�nO���j��X�(_�`��z��c���}��\K�J����ZY�V|�}��'j�{��om�9���P��i�;�2�V	l)J8y&���F��0�=zQkU��:-Ͱ&>�n�7��t��񧞅�y�2a-�%�n6�]����|�e�.�bY.dH�.���Zpω�τ��X�|.�k٠����i��쮣���gfM1��^;pn&�ΰ�3Xݗ��%j����wp5���ܭ�ly����q�a����2"Ń*1����{�U�U�n�yi����1њ�,���r�R�>�_$� H|z�� "��x���G�;����E��Ļ���;e&A��f��Ad�*�������X3����گ.�=�(� p�	�-� ߖR$.N�ڹ�H`��$ς������a�7�I�Ò}5�Ih������5�4�{e��z1��@�lS1�O]�B�w����
�B�Zc���5O!ծ(��!\����Ru&�z$0�����mH.�1�>g���!@]�|~�|M{�Ho1*��F^���-3�E�9GM&����[1�6=n��u�S��ɦ�,��_�
t�s�b߮z�,#���aĨoc����>"ypjԩ}�I��OQ~Y
�6��'��՞�!�Ջ�o:i(vL!5�2��m���Q�}�(��m�=��;d�h	�D��R��Ո�
���Zb
Z��$�CbWns��/�IP�7����\=���L;dzC�>�׸���޾����]��aJD�b�kB���D�n#����D�d��w�%5Cvo��W�o�w뫍���Ɣ�"ri�@� ��R4�e�De[1����9~;�k�9r��EU:����M��S�7O�֍+:�ʉƶ!��X6��7�1����g��A�+��ݫ�+�f&&U;0����m�xv�D�w�}_�m"BT�j�s�I�3��1~IN�ն���Lu�"N�qR�餆$�W�. �z��ם�4k��t�.���R�;4�)�g�E���ȝ]�C}��ȗh'ҤeY���"�!W�ty�s.A���Yo��z��L��&�R���ء�?�d�� Q�3F�r��Fq	�Y���/2�v�Q�|с���i��c�2�'�ҍ%uUФ~��{�Ju�����(V�n��q�lq�Xw6�?M��r^=<�����,��VaЎ{�o���_׆D��+gb��݉�xJm'��h��SUDGq�^qZ��h.��$a�͜+�Q
@�S?X��g�̵]le���ul.�>9p�4�|I퐾��-�ա�Ĩ����i�1O��6-h1 e���D�>U��ц'��EeBn����{��R|$��`�{��� 
C����^�ca.�*���!��Xi�����OF��%�j
����Yd�36������h��^���"��p}|@��=�|X�����y���Hq+��f�V�hV��-�(�o��-�	���Ϲ���\��7'*�G���^�����pd�O/�'�˹� o n��.��۳W���L�ʊ�>y�`�������[�N�ziL�q;��|_��f��[y������݄
_ɴx3��ò&��p������z��Z�=I�Y�j�?Ⱦ1O��cD�N�V&:%8��Q�xoy�#f�O�`VE��hر>�O� Q:�!��^S?�P���XߑzC�͔q��y�M�Y��au�.GC���.U����g0�f�~�%~�� 톤T���#(Q�_ÿ�[װ���lz���%��d��B����Bws*�fʰ�4�Qah���)�j�@?ˮ5��F<"���N��`�\(O��O�����)J�M��A-��l��b���ҍ!��������D5�ai�J�r�(fi���R7m�%�X�;������ww�7�Պ�.G.�+�4t�v���j��LA��������M�"ո�X�>
k�A7�z�ʾ�˵$_ή�_SS�!b2qհ}r�(���´��4eݖ]x��Lq�1�w�!�q��I�e�&O�6~#?���)��8<,�8���b\5sIK��m�a��i0�G!�� �b�Sw��-K�vC����\B�h�L<�'g#��kYN�S��4�����}ڠsϩ�5�0��3¢��C	�dք����W&;{�'��V C�m`�b3�BC[�=����WcM��*%3�GV�����r��%U�)�T�UG~x�����N���T	��j������<!��ds)����vfѠ�[�H�y�V"��ha��R͈2�k����
�&�,uR�ϟ��$�H��v�j��G6ip*t��':E"y�Rq�SSx94��bIe#�M�5Ov�;��6��s��Vi�O��Yf�f���/`S������#���j�$U �	�Ӿ�yߣ�|5��u^��H��btY��p���m��AŮ��v�T�4��_�{$C����B3(eq�w.�8/~���X�«���@ٟ�I���}�yB�X���
� ��a�Y�tG�.�������:J�(i<U,��Y}���YhUhb0��������BD�I�#?;��C�7�Y+��%�q���� ����z;�J?r"���'���]����({�v�Ʉq��P��`��_��	r	� ��񐴈��-�������F��-H��f��dhV���Ú�=�<��!�+�c�����׆���G+�x�-�gku��+N/����V��*o��j�����9j�	B`o���Kk=Ȑ��uzj&s���V��-R�F��)r�>��Ux9��q�
�x����9�s��)����/���|�ҟ<�Kjf�He�M��sV��+	�V#D�S-D
8&�G�I���-��2�J�ylI|(^F����aħW��MN�J��� ���*�ql��A��ﵕrC���m��k(#{}W�������~4'�e:	Z�p��)�����i�G���_���
H��~�����:�yO@^��ڸRH{��b�8{ �U|h���@� 3�1�Y�}t&�cDK������ſ��)�N������XPA�:����E���HM��'��>�Q�����DH`��R��%��@[���)��Q��L�L�(�q�|d`(|��%��u�&�o��j�Fa�e7~���r�v���r_��f	,c��Z��#>���m��6� ���Y���*0L�f�4��W3p��]f�	�ǚ6�E/"� ��X;f���N��4���s��\Ρ��9��~��t*e���$!QK��Ǘ���*b�s/#�`gD���ǘ-2��9��cҗ	puK�l��)V��+��h������Mg�oPn5��z�V�Ǽb���	�}J�O�M����cu��	����9g��-�Y�8� �+Ne�Ÿ�Ϭ�6��N��vÒ��T�v��b��7���y��fMw/j�1C��h�i����50�9I�T'o2�,�u�鄠�HNџb�R=>����;�m��E]���J�&�8���I-n�gɥ���O�B����@�1���I�t�e �;�u��pJ�gAx��͈�/�^D���n9;�Z���+C���I���p���{�a��u�/,� 7����[��d��c#�{9:��1�o��߽w\���'9��+��$���q�0��RKѾ�����)@��=�ph_��?�p$5��1����T�Dn�֕��B�)O��4~��{����nVw�e;�]]S p� �p��(����3�bW����d��+G���Kˣg�!I
�+�"��w����%̸d�}?�64^�m��"*��^By����'��0^15������	����]ɝ.	���'_�D"Yz��1 5{�C�Ƙe�:����G�H,�*��C��mv�<����LCHJ�LV�X�E��k�]������0��%���-���&J��U� ���1>�����A�O���UB�B_��9i����.vp��ͳhj�e�l�8.i+ʟ�����#ڲR�MW˖
�m����TYgm'�1��8�#��39��G�[��F��'�3���`W�������4.�ņ6��56Ι���`\�6���73�+�ַ���hX��%�Q���X�p�r.�ZGݯ&�;�.4/���8��l��V@��P�/!(wlJ�E�yf��W�hQw��M���L�W�o�"��_	�����1����Y3N����*�J�G��~���%LK&�|�5��&����D��Ś�����3K�V�mf�ZO$��g��N�F���{�suYĚp���$fKzN������"$x��lZh��x�C�њ���B���N���7��<��E����z�CG�Z �e��1�Yb(5�}f�&�A`�QP�,���]�6�� �2]}��X�^S�c�`����f�0�(1��������G��*�k����X`X��m� ?lWٵC��!�!n�kN���O&@d�l�)ʙS�~����U�n�wQ�ư�O@	5�+b��/�,-I��yOQ�i�vߖ��~?��$KT�UJ�!>"��̪�2Ӷ;�j�5O$-�j��L�/@;A3(�u���u\w�S��J��Uӈ�"!.�&�b)|��tL+�HqR=w���@�:�o�T��F�p�Gw& ���f�k�w,��A�;󴃿W�`#Mx�����C�������������줱���Wݑ���d�v0���"gк�����7-����Q၄r�ePj�X>b�eC��{�����m��-`Rk8Qt�^��!=����4�vT��3K�CYBg/�?H#jd�Q�_��%V��������_&���o���A��Z�d��Cn��~ك�wE���n*��D�i�Nsg�l�4x���ה ���۩��@>`R�d��f��țF��q���WxE�����4;0t��YhV�I
%�
\���Oě�J��+����+��3op����ne��'L�=6`>��*��It��Q>����W��:����^j����5�L��u�L}9:o�f��I��Y+��%IYh<�pd`��Y/<D�n:x�ު1���s�w��e��Ă�\i�<�5��XG�C�iOpJ?���3��~�B�aa��ػt��0��z�zR �b���=��X�r�qc�E������X�r�R2i�F���9.)��׻��66.܌���H�T�j>�V��=fh!Z��B`ːd����5'�y]���>t~�^뼆Qk⍦^���_�A���@�.� ������38�)ޢ�C�񍵟L��F��߲� Q�6X]�أMŜ^3{���\�ol��:
����;>A�b�^Jz���ŠJ�q;�,�̑���%U���[8�
�1F =H>��\f��0t����σ����n�tv�=@�,FI�_p�D#��F���~��S"��*�g�m��`(`������޶��R�6d' �v���!��U�m�Ȋ:�N���IU+R���paQn���<+)�J�	^(Yݥ�z&�LR���P���ȉF��5W�w'�g��\i,W�x�ZbF�7��������(?�c�G�j�]i�'C����籽7A��F�`F�d��3���oh2���W.�,��_p��v��u�oڬ`�w��`s[���`�С�?�"�$Jx��S�x��h&°5��X�`�'����8����a�CNLz�S�Wu	m{�ϟ�����$.=2���nT�0-���K�"� �!�|���"-"S�騰^��C��Z.e��l��2��:��ܨ�c!	 �!Y�~/�\�%����{w�b�M�V�o�cL\���JR���+����2:E�*�$���
�5b��T�e]sW0�^i��
~+0����XP�R�n�Q��`1>6���Y�V�P�����X�K�ts3>�N_ь��	�E����pImZ.A� e2�������XcJrF��"����j��Fs��T�Y���=#hw$��[�9���Gq༯	1�om��� `S�{go�6�@�	i�� �y�k�cK�$=
�S�����uī��r��N����Y�<�wR<�6���g��l1���P��_G���vSg�]��[jl��ؽ!��K�0����.�jUU�[-�p���DY�E����0~��ǜ��	G�{+�&y�G.�qܗ^��X�iU ?7Zwy�������6�`�t{Ђ%��?`�.V���x:ᵠV�O�"GO�O��K �V�/�W����X��>D
q�Vc�:Wc�Kᑻ4�=�lG;��k�'&���oNQY�|1 �C�bc8�1 �,;;�v_�<��`JU%�ֽ�\f�K O��	y�n��"��Z��$�r���v���eMВ���ӹHn��Eg��-#wu��q=�x��Hܟ�Id��ҳ�Ғ�`�y��1o?VQ�?�}���4�pd0�ށcv�V� $W��D���IJS$t��>:7_�Е.�p�i��Y?Su�\t�}�|���Qvlj��[_p�HO��M��J��b�Þ�R_���Q�zh�&I��6�l~kU��>�y6��A~�P�r-Y�����Ң��d��օm(�r#̟���s/������I5�y��kƮ[��5�g��`>�'�f��E�H�񱝬�&��@���d���%�d�Q�}����(��$Z�S�j작og��Gzf����ގ7�Yk8(�pܼw�;�	�D�_�i�q�඿��>�ه�1S{�����r�Gb�&q&�O��*��M#G��+{p/�Z�����6o+Z\3h�	�!��h��:=�҆#k�<���������'�`o�s�fZ��s�|W �R7�t�iӈ�C�{ia��\��X���B�[3W�!�1Kȓ������=��(!���h^Ql�Tgc�V�����'��!r}��w��|��������-�d��SRK�R�$���ֲ"�?0�%# ��s�JA�qQ��M�Fc��~_7�p�sAW���Bt���]g�����|O7'Y�hH��:T�p�4���	���ܠ)`�ۜ����W糿u��z�dٌ"���P81��ٛ<9��b��3I��-�b7�[�-�TD�	�t��6@�b���$ �[EO�FFF� T�@��˷:�Ե�k�����LO�ʈ'��\9^I�l9͙ǸPF�i+�@���6\:Ma��f9�1}��Q�#���	 ��(j����7
�Ӛ��R��5��m��CWK��-�=�A�pD�Y�K�nTpf1fȔ�0���O�j��G*�?f�d�w�����i�uiF�p��D��U(|�tɋ���`�ץz��ķP��<�,n�zAD�0B*O\��R�Wd�Ǝޅ�^}������=᧾o����Έ�܈C�ZO�A�b���EC	����>J���b O�E�.����`:���q|d�Gp��_�(P�����Cɲ0��.��2ﲁ�z�͟F��I *��2��=q>Ls
4�&HĬ1���WF��t=�c���0B�~w�6�*�i@�G�{�2�8�?(X��!c�yD�LH���]4a��z۳gLtFm:�2�N'���]�b"!G���xN�"�DW�x��k�E��N���KL6?߰J����X5��B�Βs�J|p(�*���`�븳�A�v'M�M�]�=�!�/���Y_�(k�y�\�w6�*eu�%��%��蘱�]��[/d��RoKQ��+/�Y$�͇�&K�k�f�-�{l zo�I����!����; �	��B��Q���u�wn�7n�j�k%2����d1�T
�'�<${�y��ԎlOY��K	���8�9����.�l����hs��9�&�ʾ�QQA{�ci�_�+���[�^+���c��q��>�����5�$�+�'#�_@ӂ1DZ�ک�܅��j��SP��1T/�i�sO#�: �cW_�<��g�w3Ue#�Ė#��=<�ŝ�Aq��w���DU�}���%G�k�J���=�4Q��c� ,cq@uy	3��,����q������ѴMdӝ���x��-R�)�:j�(#�l�/|^a
���ֹ�U?�t%��[�^�(�;t�gSxP\�OHc�̎���6(G���݄��}�|�fmVYށ���@y�Q���N �DӰ����P_kR.����J@?J�4 �V-
0*oO�8�VO�D��#��� W����6��h��7������}v�#��:7�N�xK-K�K]}���~�I�}�t�;�h١ˡ�@��9kyp�����;f�� �מ9:-��v��$.r@�`xR�V$�;/�=�sM���X�9j �+|�o��Y����B�����:{W�������_����3j��]�����7�>�m�/G/M�1��qgW(&#?�j�I����¶Ш�5w
�ɍd�!�/v�n[�9�!}?3��R����~~����k��-���~k	�a(-Ϥڵ�%�w��Fm�n�\��$�l"~�����l�U�N~�9�*�O��o;�oҵ��S���Is�
7��r��K�։�ZG���Vg[��\�M��{�f��=�v�ߩ1�TWQ��ޜe^?T��4r��q�Ώ�\�8@ =���.w.�\<�L�0�F"���[�%-�OKبj��Je�tt1(�J@��BM���IZ"�T�zϏ����y�u�1�Z<���~8�M:��.��u�b�!�]|\����R�"�(Gq����>>L@e�^Bu-^6afJSP���xNT<�(fV�{��0pcʝk�܌'�$E�z�(�YNk�Ja������L})����Z�^�^0]=F���۱i��8�~�y|ur�bj������&)��t.~1}N�Y��������� ��԰)�o�. ԔWE&��Gk �פ�C�o�[��4ט�繾�rs����5�%�U7�#�H���[8��)�׫�y��h84�d��ߩ#�q��* �?H�1��ൿ���MU��
�0Wu�'`�2G��-��OR��Ժ�6�:�اX�r��?B���Q8*��f/��Ps�є]4�=�E�t�������h�x����*��ɅW��a�D�q~JYL�6����X�A��rom�����������n8�be��⁊T���TJ�{C��{�vke��F��^K�����`��eama���@'�P�Y��{\�&0,�YǄ0�h��.ۥ$K��~���!�B��	���[#.�E���9��tNb=)�czD����M%�v�*���3��N�0�(r�[b,�9�aq]���e�ޒU��-��/ONR3�Z�K3N�*�=��8����J���������ܱ(��[�K���C�uy�qh���U�VoM�5FiY�76���x�� c��.��P��;�i6V�2�R˯k�����p�v�q�ɺ��Dߍ�bb�˨�ߑ@�����y� �J��P�W����v��X���8-�����g\��������Rw)�*���Ƥ�]+�$#�z��3`
�[c��4���.���(M|,��������<��)�0+��Y�c�jԋ���(g�F�"
##&)%*�?9�iЛ��=���֦{Iq4�^5z=Y��2���~��v8  ���K���غ�\h�2�]IE�s�iuQ2G��[�kO�i�X���:+ֳ��J��]k�-b>�d'r���9�u,-օ~�����v��/~�#���U�Pe=ױ��\6��
9YJ'*sq�qzE����A�����*�O
1?��Ge3�F��Mf�� lI+T��ꭳԤ�H�sz�e��[�������X욉��67<]2D�����C�-Y㣨�~�ʄ���Y�j5���S�$��jك����W��ݳ�ܽ��~��%;Ԋ��.]ƙ�f�D6�� .��kmQ̨=�4�E�Ǿ)���Ɍ&����/�"!�E����[�=��S�0���y�#w�1�Թ�l*���16]҉��������.gR;ϞE�d�i����W��0lژ;]����
.+]7�ye
'��e��ƖO��e����,E�Їe#q�2#r'I.�枱 6����g��T�8߇��um���ߒm��|Q��a�0�DE(u,��^�,�6n<��k�{>��F6�B%^V�E:J�ok���}̖����Κ	�bqL�P�"cP�-������\C:��dj�Lxp��$���o��4+cI���"9\�c�-����K��E�w�3t�zT���0�ġ�֔����UĹ�Yx��Z�+8� K-�s�I�q+f�3y�Ix����Ǯd{|"�!�����a;��x��H����׬U������0�T|E=W�0FxĶ4{1N����oJ��0Qf�?��r��q(�l& l�À�/��O<u�
۸��9I�)Zo�����hJb���~!s���|����{��urV��_&�$M�
hz��8���&$�_ó6���������Ƀ��l�'�G3߃�_[.��N��j�F��i_��7MD�Ϟ��#d�9%\�4�O��%��߼7��b������I��R_�?0�a��I���m+<Z4y��������B��μ�1͹�+̷��\��C�U��t��&�:��5�:����4�>�R��_�mj Z�X���4��d�Yɼ�H�+P����Rյ��@����L�P}覵�D۰u*Z������z�0��\Ѧ�JL�DeZ^�h��5ۮ���|��o�bY�̉m[��
�`��N�C>�}��C͚�ŠYTm�&ď�&���g?��m*{�t��#m�jQxD�"��V�1�X�H6pu~/��L����E�E�+��u$B�\6䡗�)�Y0��)�i�\�d����ؘ%6��y�76�S�[F����#�4M�Tڍ.��hB�E�%�������(��DE��]�&p<cy�e*�6��'����No0�&�QOw�29��5��
 k���m��TС��a���}XPl��'���,gB����4m�r^�{)~��n�U�<X�]�eC���m3�����N�G��N �-���Snw�a��-FQ�`w�0 v�(��N1�/�c�>��%���`�7X� ��1��;Uvª�}j�dk�ew�&�.R����q�mU8��?D�Ӄ�@��xE�w����Թ�y:2���GJ.�+���F&*�[�4Q#�Q`�
@G�i���ԇ�т�`0���c�`�>;XGS�ö�҃��ǣeSG!��̿K�1�;�Cj	g�:���󍜹�H��Ŋ�AC)d:�L|r�FY���C0���WM��(��7��r��vsi
�8��0z>݂Դ&��
������N�dE1�i;��vFp<(�B�<������g_��I��YP.2���ҽo�;"������:Ŭ�Ւ�q�4�ڜ����\����S��k< םK͔�v|lO]=:k4���y~(��n" ܝᙱ�jWKa�x����bt�$�U���jK��+,=��o��9�A���6����a=.f�Z��L����ҹ��L��Ey���Bǿ������z��M�H�XL���'�����D�8� �k�eH\h��/yW��0S
3�2���Lx۫�#9������l�6�h1�n]�����n�:�'�6\@'�N�q���UZ�1��䛬g�ʿ��BE :!�5�A<�3�2\`����������:�ˤ���D���	~�N�Z��)kA�r\��z-��@ʲL�S�����M��#)Cf*d(��ܩ��h�HS��~�� �GM
�F�*6ty$�YY0O����M�m7y���0<ͬ��%C[�� �� ԯ���}"�E��`?�K���%�\���Y3wq��"+)jח#[�34VtՇ\3{��|m|���4?�¢���(]5'�C;i����ȗv�[���Yz�G��/^[V��*�RM	�4���`T��������E�%�gƖE�g$A�ʃ���:�;C��$Q����BԵ�xH�/�v�ߤA���[�ӻ�Jf�i)t�o�o�!����
��!���#�Ш"���'
���b�Q��|l4�P�1���/�`�<4��n���z�;d�
���6����ū��ժ�i�@��)Q�QȬ���R��|0�p��d�ѭ�,}U{C�����q����e�;�qr��B\�"l���ކ��� ��&��c|�S��À%�!oԕ/�9-��Ǳ�A��щXpUN�S�f��?R��r�X'褨q���`ܳ{���$`�kH%�-�<�H�y�A4��؏=�P�E.SG��la�]��j�i��p�-{�������2�X����1�7W�6X�%2P�%u5�qJI8���i�_�lg�2�T'��62ir"%O?�x��S�9%�0��*}hRm��n)���9ʹޜV��Ts[����A�`�!�b���f���ު�N���6�md�9埛Zi�{#�B�~Tr�q�Y~�.��*�N�����(}ͧC�Q�f�8���,����\�$FTŇz��)�J���@�$R�!F�]o����9�g���4:eJ�k��[��27ǝ�_M����ܗ���3S	!�T��Z�H�k��N����Tl�c�H�	�w�ۀ��s�_��*��E�����o�{�Λ�5���熚�DT8���z���&�D�&6��m#�Haѳ���!M�zA�LH�v��%�/�*D�@p���ջwk!����ĸ;W,<���X}>��E���m�]C�!B��aֳn
�CQ�K
T�g˵$�|��F} *�Ūd�Ryݪ���}�������u�9�S�m���J38��2����G��aà��@#�Z�����} �&R8}�s��+i�\����<u�>2�.Y�"{!_G�؅���̧�TJ�q�G5{��؀���+L�r�A����'��b}:��T*ÜG�T(�a3�R?�6�]���g��ǡ6YZg�i��B�ET�G�#��8�T���5h����(x|J hͲ�0����B�(�'cK�yh���Y:��CN�o���g�̮,��4 ����K�1ƻ�x�ʐD���='Q��}˳����&ߪ�ʁo�*��)��r���`�%{�~�۶�L�_�Nt6�^�{ dQV��=n�VڕP��QE�8����'d*�P�"���If�g�����%.Ű�" Z�]Y���AG�z����p��x�1�/DjCR���v�I:p�S��4^�X��+���N0�Z��o��1<�:�58���O�[#�u������@T��gz��G��-{|�ѐ<A{����K���/-�oa��̯Xw�$R���ہ1W0l�q���=O��D��g]I�F=�����t��a.pk�Y���X"�~Ҏ���#m��{*D��_42w�����[F�1������)|���',���]�:�^���|�k���'+mW�Ш�@7�<?��#v0��Ih����r������>ðy5���~�-K<~���ɝ��QHG/�X>@��a�˒b�Rq���z�KCP��.��!� ���,��+�����[���!�t����f4>,+ɵt�Rq��Lf1�ro�N+�
	Z$9an8&��lEiM��p�щ��Na6���p�`8nz�_\�t�fp��3]�f��������"�Z"�k�Đq~�Џz<��u!zg_r�C"��	�
��wC��T�6��Ŕ��
�7�b�&o �}��SW���`����Cߛ߀}��I��D��!%��T9�a�����-�S�D]��:q�g@�P��J8,}���P�mt�\��b��Jm���`iH⋒Z͔��@���R	z>?y$s �� �A�Xr��6� �q��Y��O�R�r��?å!�R���b�}��,��SQ�gM=�g�N�c4�z�I�%�m9���F��1�e�i��m��/��"���1�t��H�fe��^�ٝ��e������5E͇S����z�Bl�P�� i�a�K,UcF��ق��#���nN�����kF��46�˖)�wbJ��H#�p�����{2qf�ݚ��e��ouiM�q&�7:�]!7�y��t����C����EL�� ��S�#=GRA�+s��p���*�v���o��)vi#��>,�6B*\�kk�&r��Y�/�RAM��>����~dlX��k�y�P#8xEdӺ��\��g�`�,6	Q�_�
�	Uɣ2	l�/�Ф��g�1~�nd�iMC4X���#��x�C�q ��,����֌�Ý˸�@K���O(7 ��HC���ir�AU�ތ3�?��;a�:��?���E���+�r��\9_�����)\�5�f8k"A<��.c��+ă�O�0�,p�x�����MB^����@��	S'��J���<�52X��ER@�����V��������J&�!����ᶛ��X)oM�ۀ��$�C�I�]��}w�Z��iY�Gm�%~jݭk�Nm�v>��V�g�Fq�B�O�N����,W��`�D=����_m���u]���2�D_�Hk��k��6g��E$�[�Yd�vmzw�H�~w9��9�r��xD	KL����J�	=B(�,�J����Ԁ���;�Lrl�4����>P��L�c�����ԙ,��@���zb�|��~�ѸWAo�E���Ы�W����)��\����%`�ˌ}���~9��]�N�(�d1�G��ye�T���DU�
%KD�wY1y)�)ĳ�/X�P~8�	�>�j�Eo�ܦ�:��_P��K�Vs�,��h$��a�e��]n��N���`M�i��[��2������M{'�~��c��2���:��D�:v���tM�G���\1ď�U�(Y���ߝpg�"�%�;�ڹ�6����oHtD$|g�A�"(BM:��K�a`�*o���,#�����A)�!&K�&9��}�<�`�Gۺ�^�3�#��Xnd�l��*đ��t���İ�.��O ���C���6,��X�A�Z��z˧1]Xg�j�T��@�8�?w=����Aƣ�ݱɅ_���������ȡ-E}>��	�(����<���������<���2���a+�t�+�3��)\����2@���gXQ["\�C*@��\�`�G��2^c���Y���]W�����d��
�:1�����}-a��4���p����CS@&P�8��M�vXDW"@x���=�*��(k2CY�˒�F�}�:F�y.8�p��Wm�[���ܵx��D�]�N�
���6�V��5l]-�/�g�v`�!]��)����Մ��D��{dRdv�Z����)-4�o�`��ҝLS}|ݱ��_��(��p�����޶O����|�Q��FV�/�t����G����G.F��e�}g��ۨǀl�ר2�$���g�e� H���o%����&�� ��L���_a[?��y�,�bt; a_�W:	�X��͊`���4���6�C�<VB�H��b��O�|��6�.�j~v_װ;8v`�DL4W�B>{�9�P�I�8�n� Qr���wƩ8�������-�ۧA�M{z��V>�uv�5��*������I�������л�����P�3��z4�qa�s:�e`ԟ�DX�3t��)� �]�yR\p��o��͉��Dc��G�Fu#�ʅ�h��3�&��0Z����w��¯�y6z�KS��
���ӈXU�_��JXƧ�VSГ�K��K��y�[�E��~�0?;��m��f�s)��q;���[F��KK֪�.���+}~<	�/�_�l, ��FS�T2��)��Mp4����3�*�6�@�u��L�l╌�4b98�;��������	�8�'�p0�[)��!:�p���H-���3�y�:�� ���Ђ����������}G��NI��(�$�oj<�f6-b��Mhcv�������v�P<�PÅ�/᱄I) ��ϐ��I�x���_��͡�}���ڙ�"��g���r�2?���6�A��R�<(w�fޚ�Ql��ʽ���Z�x�����\��6����fx�