# ====================================================================
#
#      altera_avalon_28f256p30t.cdl
#
#      Configuration data for the SOPC builder aware AM29LV065D flash
#      driver.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####

cdl_package CYGPKG_ALTERA_AVALON_28F256P30T_FLASH {
    display       "Altera Avalon 28F256P30T FLASH memory support. It can be part of stacked memory."

    parent        CYGPKG_IO_FLASH
    active_if     CYGPKG_IO_FLASH
    active_if     {!CYGHWR_DETECTED_SOPC_DEVICES || is_substr (CYGHWR_DETECTED_SOPC_DEVICE_LIST, " altera_avalon_cfi_flash ")}


    requires      CYGPKG_DEVS_FLASH_STRATA_V2
    implements    CYGHWR_IO_FLASH_BLOCK_LOCKING

    description   "
           This option enables the 28F256P30T driver "

    compile  -library=libextras.a altera_avalon_28f256p30t.c

    cdl_option ALTERA_AVALON_28F256P30T_FLASH_DEV {
        display       "flash device"
        flavor        data
        default_value { "default" }
        description   "
           The name of the SOPC builder device connected to the flash 
           driver. If this is set to 'default' 
           then the first device found will be used."
    }
}
