# ====================================================================
#
#      altera_avalon_uart_comm.cdl
#
#      Configuration file for the Altera Avalon UART comm driver.
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####

cdl_package CYGPKG_ALTERA_AVALON_UART_COMM {
    display       "Altera Avalon UART comm driver"

    parent        CYGPKG_HAL_SOPC
    active_if     {!CYGHWR_DETECTED_SOPC_DEVICES || is_substr (CYGHWR_DETECTED_SOPC_DEVICE_LIST, " altera_avalon_uart ") || is_substr (CYGHWR_DETECTED_SOPC_DEVICE_LIST, " fifoed_avalon_uart ")}

    description   "
        This option enables the comm driver for the
        Altera Avalon UART. This allows the device to be used for debug and
        console input/output."

    compile       altera_avalon_uart_comm.c 
    compile -library=libextras.a altera_avalon_uart_init.cxx

    cdl_option CYGPKG_ALTERA_AVALON_UART_COMM_CFLAGS_ADD {
        display       "Additional compiler flags"
        flavor        data
        no_define
        default_value { "-I`cygpath -u $$QUARTUS_ROOTDIR`/../ip/altera/sopc_builder_ip/altera_avalon_uart/inc -I$(PREFIX)/include/cyg/hal" }
        description   "
            This option modifies the set of compiler flags for
            building the Altera Avalon UART comm driver.
            These flags are used in addition
            to the set of global flags."
    }

    cdl_option CYGPKG_ALTERA_AVALON_UART_COMM_CFLAGS_REMOVE {
        display       "Suppressed compiler flags"
        flavor        data
        no_define
        default_value { "" }
        description   "
            This option modifies the set of compiler flags for
            building the Altera Avalon UART comm driver. These flags are removed from
            the set of global flags if present."
    }
}
