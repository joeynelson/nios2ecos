��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_���Ч�;.������1q�m�˼�Z��6�E��H��!�)�-��*S=����C\����z�WOtj��4	:�x�
N��<��K�����N�J���+[�S�ߊ����J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��W�Q��L�Uт�X"��ؖ��1�O[�B���:��B�X]U%�n�g��5����͉�׃PuO�]��p�>6BD�d����MNM�è�%���*Mw��s?v5��P���]�]�$������[�>.��a��B,�g��Lð�p���f[����R��ix�b��B�?�o�r�hV��L^GR��zҀ�C揻r�K�\�>����q)u͞����m&�(��G�FY=�����ߝ�@�b`�*�{`�3�n ��K�31���G�g�r�1�Gvd{�t+C�X�J��\P뙏�lBO��9�����s`���e��q�h��c�?*y˨���HI��h�>��R?e�YExgU!�Z�C�>!�S����R�Vȼ��K�V�=<��A��%��[8ʔe���k��*H��ej�h���X�R�n�DY�%�zp]\�:]7����D5��K�2�nWl���zf�����*�9�K�� �Jv����`�A8,�ڂN"�E�� q��<�ɭ��"a�Wx�/�~��h��V��<Մ&֊*���/ w����c�
����p�C���37~�DvQ��vh��(Y,1M:b��8��t(�E�C1K��a��&���L~R4,�|����z>'�Z�p�{o�=�kfE�N�3J�<���&:x�i.�UY�Y������� ��I��ε?�9���y7���Ht�w@�tfiǸ�Wm�����B������5,��	M�%�J�)i�͎@W�N�`��S�˜�k9 #��R��(m�n7b:����Z��Ά��ƽ��٤Y*"�5��Q�s�7�:�[�(��-����ȓ�z�鱼}��r=��I>N�T\[r&�	��Ţ���%Gkp��d�Z�bV�
�`�����"�i6�z���KC}(EG#C���O3e���Ys
�rh��5&W� h��a�l^&Y��H�8�j;�lv|Z���Ҵ���Xǻ���x��GUy��9T1D�W�Fl~@�:�%2���6�g̕�cZ��9���;�(Җ��G)�3y�N��J7�Gm�Y����4X�� ڻk=�M���j��#2U�,�Y��.Ĩ���[�)����;�K�T��X����c�W�~H�j�:4�&·�����d�s�<�?��tI]�;�}`ڦ�%�(�C��X��>'~h�'ė�^D�'�`�'�t��@!��ʞ�n��z>��cӑ�-�tb�4���Tv<���v*l��h�L>i|-Y��[����a7l�2�;K`��f���L����x&ٯn	&.W�D\4tr�u!}|�0"��2�\�;��� ��ٶ�"�]�\��Y��!a�/�r�Er����a�<���gh!\���uI(/��W ����W��o�[Ґ.kE==Ob�0���;�����R���&-����/����K9�@T�߽I�.�w�����di|�Ԛ��ׄ;r�d8�u�8!�.P ��q"�n�˟�g��M�e��E�wf�#�v�a)�"���7o?`���6�V�]]����M���gd	��{t�Ӝ���1�n��}�98�=���|&�b'<�έ����%?»L�}�k�����'���x59eS�h��rR��^�r:�K]�Jh�u�4���	VYA�T�roϿ"�0E��%�/��a/�qk1U�Cwj}�xk�N5Qhj��{��k8�|�Yqv*��d���j 2�	"f�6,`��?b�Z!��M�;�uR[�U���a�w9L�,Q�t�,���0^w��#W��վ�\�dNl����L�[\�-a�,��?>��@��-:s�B��7�#�����s������Q�����P���E��_������DI�f���9e��3����lo��9��݈�������)��I�X�E7NI��u�u
[<��ߥ�6�
g�%�l~�Z��.��N|�Ci��� �|bF���Q
��y��,^����VU�As�F�h�m��E�LG��zO�ȭ<���i�� �@Z�Zx՜c� ]0y8"j>n��p�ɟͳ�zW�l�݄�1���T��8"ő�h�k#Eo����Ve%��p6����ٜ[��s��F�7-��_3�����_�%���_S���F�nv ����}�@@�6�hK�ׁ`��������Z+J���,J�粀ᑥ��V�ݳ�X���B`Z��G�~]����2C�Y3���P�
DW�߲E�7���gf�����E~ɞ����Z��<o�4�j� tͬ�Ng�7�����OBW��[�c:���w`x�$��M��1���ߛcf��N"�?�8'��I9@���3�����f�M~�Ձ���r��N<�H�'��G��-��"��oLK���� ��)��kry��LB-�P�`v�b����>] |2YlBs31�u���Ej=pA�O�}֑j�2�B �Y ���u�8�Ƌ��M)�Lv������K4Uv��h��R3}��V�G2�����F�ʵ��Rf��o�D|\������ǣ+-�8�"�V�2�e1bW��ۼ�|�P,F�/��
f���b�����D�т��si�q�/U�Zlbʊ�A�G.P��8$��rk	~���}om+rL�*������Ԭ� z6���b�ߓ�����P���G#1 �;��Vھ�,�3�!�If�t͚u��Z�)�n��~�����5�T��Ͷ#���.��c��=�]qν����OHb�����m#=��v,ǰ�2%l��X�'Qj��|�7<,"h�G�P�
��K���v<��׎_�^;�r�֢����^l�D���f��%�1	.������љ:�K������Ꞻg�1Ȅ��W�\r޲��F��00T��|]�/�0~4h�C��VQ�Ʋ�k��(����N�?g���|��� �M�z&��r�5��%؊ƫ��-��v�*,,�S@�A>������݌���>y4=|&�ADЇeB�
R��Mj��:�$��؝h�����Crg�ΛM����_T%_�����6��P�ގ囔D�Vi֡Rdq��΢�=`7����'u|kW� ��x��X��S�X��ÔUt�U|���\�P.`d����â	K�{�!��ܝ��p�=�-V]�dU�^����$SG�ܥbƕ.���/�g���j��3c�(T������V�n_�Z��&���}|�H\��=�T��:q�0�I��*a,o�� ���� ��"a��L����"�G���bA��پ@O,F�h�W�V�Ln=�������fH �'��C3��g�ˡ䞥���xfK�VR�q��b:�e+4.���n�o ��J)���cC��i�5(�m �Ќ����9���45���z1\�hELIU�+ó�l��J-�����¬��A2g�(��Br�L�n��"��c��t��x�z�;��(8������q8�˖5]n7~�
�n����e��ըO�k�NlE�hSUa��6H�t�iFۂ�2�(8U��lM�ʩ>+2�?�x����W�m�^c�x�A�2�^���b	��B���Q��w_�"����qs�,��L(��t����݉R-T���|V(C�"G�����d���r�Q�4�mk.��>P!�uzG f��zi�\T����$y��bE�����Zi�>��y�j	c<Q��T�|�(A��ֳ�V�덃L]@�jԷԿ֍v��䥖�@.b�2�q�Zq�M0E�H������9{�c�R�ZE!ؠr�w-e��� l�?��Cv���ӑ��1��� ���_�Ȍ��[f��/��Ox:�
^?�E�j��}���wswq8��:�9�7�ov4�>�ig�u�TЉ�Oa����E9|1QDQ_<�R!��.��b���m�]j_>�����.B���b���_�nI���<Wd��#ݭ|�wS��à<����2�w��V@G/=��(k�H�?���ΖI���8��i���7bdʗ�I�����J��e�́L�3hR�G���㌞�?��a�!X({��
� E��GH*��w����rxk�j�;r��u� ԿTtv%�QJ�ث���Ӄ���$y����h X�o:�^�Cۚ�4)�FDK�~9rl!�6�0�5��ϟQ@�jZ����wv�=����4�w�`.��Lyl@*�䝔GOKX ��ݛu�S�K�qw�,7	�0ڨ]�+�tce��"|%B�}G"-ck)w~D���������(y��X�jc��
��-�����h��E�Kc&���28���*�y\I�H�v�O/����M�Ic%0�S0py硺��̊�^�yiƸ}c��\�{ܟ}��0MF41�[�kJka�Ɛ=�
�&*ڿt�v#c�n��?Q�H��W�Z�jfC��a ��f��}���ih
4�IWa$V�&�ڡ�f��f]��!zS\ 1	m>@p��ni�.��0?�}�k�k��D�ϋ��o	��fml��IkC	d��hG޷�x�p��ô�zY�U�J��p�ΊGo�춛�#��k�
DQ���P�K�i<<���c}��8o��s{��7gY�%6�t��/߁�?��Y$��8�*o_O$<��Ò]�4r���D;w�#ϊJ( pj�]Y&���~t��X���M���r�Dȧ���h�ԏ���܄vp�T���=[��:��n�:�ǲ��*"����Y�Yb�*Ǟ7K(��)�L��| �����S*�!�8G��,�G���E������ogxzT��;}������B�Hd�R�?��2X�H���w+(����,�4U6��\��+��-*�#�8�ֹ��tk�����Z�-�z�E�e{����s:�[<��óm�Ȉ��_�L���Ţp)����+(ҫ��/�����_º�d�&�-�oY��!�3:��k�Pv�K�]�^Y���n���ao)f�������	&N��B������:�7�S����ߥ\p�����d1��A
SH��bS��WC���4.�#��A>:ɑ�����9c�EE�u}�= Sh$��Bt�Wv�
�~,T1��*��5���K�����t�ۂN��ml�ܦ���x��1�Z�]EB�1��8HZ�R����j�S�gs����@?���j*��x�$O苋c�M�h,���N�(^�b"��!HUPo���::c���|�Z}Kh /&�=qm�F���U� 2a9)C@�~��#.�� ����Ztt���z�aϾ�z�3���������Nw4֩�������n)�r�G<@��Df��׾2�,`�{�i/y�-�[A�/��XX��WO����fl@URf�j�����QW�M^<��4l�Pw"�.Mo5 �(@K��5��ŧ�T�YR@}���ѡ7�s�2`�֪%����c���ڣ��Fg�|7f�l�|�c� r����Z�_%�ݜɗ�q�X	��A�����M"#�������R���I�i�E���e;�Q���qjs�yC�.*@�����x�,.�?o?1�P˝�,����294�D�w�LEb�!OT�.!f�:�]]�Ӿ��e]��&-�r���gZ8f�O nZ�E��jxk�aI ���7gW%6��GC��>�ܰ��/�V ��ML=R�@r�_G�t�k5�5�z��y�E�Q2C"���uC������luJ=�Ҥݭ�/.v*Jk��S jN�U��p`�v��������6�%�:C�P������$�t����-T�K{�\�uA?|�̼0s)ť�;5�{�:�}?PP��Gn�"9�g���F�Xh.��>����02Ь����6��;�΅���H��B��uz$����FI�Y����u�2[��e0u���<�O]�D��_W;�q����b&�ϕ#��,�9KP�Z�����]e*�yT�J`.A��}C|4��	�o��/o:܌P�PVZ�q^��7�rF�'P R�3x����D�����Ƣ�M��eGi?93t�}� ,{��	�i�*[p��W)�'�H߲X�����lwo1�f��gt���D�!�$��#bɤ��Z�Rou�+�2��ϱ쀘X�����a����m�]��܍Q�)�o���k1�~-�j�O'P-߾lS�ov ,�3ʷ*�6=8v�G8��',��j�喇�2��0Ep�?:��QI-
��l���	�.C�,��
�V#{�wa�4X�Vj��ڔ��p�z��ޕ�.hD��Z� �cV���,���3�^�]o*�u-������<�w	(�^�嵷�ͯ�r+e/�LM/?��1!�FZ�۶E�&o�,�s��+�,BX�ɸ�>�$�$0������e��ms����D�4��xm!j�llD���4Z��$�C�]�*���h涰��e�/��u��&�$�ϤF���0R�̴q���D٘����*7��BY�?�I(�7�ڽ�����X�j?1�V*��qި�e��"�#!��m�6$eJ����5��k /J*E��ߪ���ۢ���e�5/����r���[�&*�������cBX�A�������&_�E�*�r��I����؍��G��V��ִ\|��\���6�O���N�;:��b�ML��Hz�E�Hw�m�G��f@f�6�(ԇ/4�ڠֲ% �����ltR9q��HK��u�#�B)���d�GY�<�x��O�
7�f���9J<����"ί���#;��]x�K�1#xT�I�T���9z��Z�3���OכFٶ�6��dߦ��z�L�[�U�$���M{Wɩxf�iQ���F!4�:Jw-�HR�pW������
&,�N?o��F�bJzS���p��W,���/t�{�(�p�զ���T������BW�t��!����F�i?�&��p��Y�1��\���!'q�z���g�&uĀ�%!��&�ad�*Ɨ=L|�vfJ(3@�V3��`y�c"�'P�r��$J\��\�ݺ���P3�N�q��ngrڗڳt� @�H�����_�,����k�5���#@.��Ho�Ρ{* ��x��$�2�_�
�<]�����=���G� p�;-�^��D�b�+
�$)I
���D��+�%�y���8�'�����+�����f�KO[��p='��a�;^F�vG zYx �#L>�����Y?�5R��dP��G'3�Q߅�Uᴿ]A�,v\O�/MOSq�KI2sj~�_���	�x�Ѷ��W��DX��ojqrz������K�Ч�E��0�����~ܽ����F�LU�M�M��n��>���R�{/uE�/��9l��_��������a���I"9Q�Ey����|��Hl|�����ӨU����.��:�+	n�p���D@_B�t(JF֊q�k���s��8�ɽ㰁F��Ce�t'��y�4Q���8�ߨk:;5��M��5�}NxD���������F{2����hEt�����/��Մɡ
�n��_���3�ׅ���ɑY\'�b��K�W�gw\�씝�^�Н��A�u���WH���]�ҡl<�a+�^(�;%������Є��=���K��<|�v�,b���D`��b�!#^��Gb(8����w"������s �5�K\�X��5�l}�k9�ɇ*�s��:��$��O�ײ�x]ڥ@�n$a�s��(��M~�q�<]�e|��	w�:Y��uR���Xۋ!}(�s2g��O��WJmF�nH��e���f�h
��N�ڣ�:�_:s�ʎ�_�U^�2��"�@�Au��70��A����iY��˛m����or���,�G�s�~����	�:F�*��&}�e =R8��DPX�C9�[�=��vp�
�O4�5H��"�X&T��-�3Z�挌Ҫ�Q�_��Ex�-�8�a�n�0�V��f�:D��L����HG#�?<R�5A�<��hO��:�=^�8�.�����Q�pѭ�G~�H[;����N'+mAwA%�6���G���!�d�Er���#	¢�_d���Ƙ6��������Wu:�!���-�9� -���| w��X��|&A�.J6T�։�,H�»��b�����a�h�n�;�o���M�T���n:z_3 ����e�X6�e��r��`^P9ZP����˼��#R\9��;�.X�3A��Zkh�/�B�ks��� Ou���C�P��p�]�¤�b���$� \��*�s��/�|F��^��d�D8ւ��u��8V$����u���t�J�1��g雅s�/)k;�Y��[���ڮ�3R�t/�Y��`��"$���0j�'7��i��$�o;"0��X��y��)�q�'��=�̝yo*W/1�3��)f��:��p?�j{#��ory$o	x����״���@]<;F�7���zbU7�=��ȩHkx��Niw��ޅ�BJ���\!m1���� ��A}�m�%�#Em
��YR����׳&\ǂ�?(p�zIatn#8&�Pm^)��TB��}�Y�r��ً[�=�K���� S��'�"����L~����L�Oq�tQ`|�%6�o�Bqǹ�<�b��_RPƨ'����Q�����S�C�\q�i��׫\ur�+�i*����נ���$�g�	�m�>b)���C�g����:B1�M���h6������_˘LJ:L�2z0a�i��lOR�+��h�*�e;1�CS�n=����!���ꗁ�=u����Y�K}ۭH(��'Q�~}(�b���c��L�l~�"D�����_-ݲ'8�<krR��D�SL��0M$g�w�0�y�[W��B� �l��l�b[L�F���2z%܌Dϳ��!�A��.�N�~��F��ux��>���y�d���F����	��R��A[�42�
%	���|ez�J΍g���f�$:��!�`5����#�����lOz�`r��lQ�TY���xI4Ta?��	nͶ8��)4_SUTI4��f�1�/��x��a�J*�zSǂZr��Ҥ��%E����(u­6Ex�Wj�\��}��zsoqT{��믈'�=�
�ӓ����F�M��h $�0|o'�� *���X+��]Y>� 	_y@��������(�X���w����gCZ��A�7怽I����W]���*ݕ�����xQX]-�g�Q��(�#ڕN���7��|�&���������i�ɻ�U�J$V��7�E����3���\�ї��ug��<�&~��	��āaQ�!Z��[]}�mc��B�e;��@�Y� �~	��F9��N�g���#�a��7h >���秢q�;1�^)ic���s���c\n��o(�����i�۲`s�@v��+:����8��}x���0�v2�_Df@��k�Cq Ԧ��V�W|د_B	pJZr��>tq��Q_I�k��A��<\Q1�J��c��Z4y�:T��ro������:R���}�ϾG�@�C:i'�(������b����p�j:�A a���K���X�+b�K�E��"V�r�u�}?\Y�Dv_�~"��6�����I�A>F@� �b~�ȌMP��a"1�B��d C
��Ac�6>� ˋ�ڝi���k��9-�.��ۧ�˸c#�w+�}:;�-�D���+��\ !h��4��T�6�GFPV�ag�]�~W.>����O��C��8�Sm��g�|�ץ<�����B���"
�����eGA�.��Mcm.؈p2�6:5[mma�w�;�R�J�:�ä�|�%��qg}�N�Na�A(��(�9�~s��t<tV
�o�-�<�7��$��Ԓ�0�:���7����H�d����1ʠS0�=>�kۅR��:"�XO�H��B�c�ũ�ZZ���MYŶ�}�OmH$}ӆ�g�R�9�y��ew����wm�ݢ���ȳ.�(_=��\j�`&��:EQbģ�eQ	F�Q#ͺHi6N�,L5�̴�����S�N�tϖU��C�e�����d.O	���@���6�Bː�#+5� wJo�]Pn-��	��)�Xe��_^�F��ɬ�uvd�\�ܙ�S���e�v�W��A��a7 Mm
�Dvx�6���H�ker��5�rrf
w���>7���p��}���%.�&��hY�yE��,�X7��Qڎ��F \��8��t}#�{w0Y:L��Pt�L݉"���d��	@�8����j�rBA[D2g��@���UN� u�����$a jQ�)_��/}�>������o-��6��Y���	�z|���O��I=���� ?�bnV�t���U�2Ubr��Th{�g��A�@�}�(�J�x��҃�:=�R�-�˓��W���� ���S�+�#ۂ��Bl�����A],�ON�E�n�i��`�	�ַ�߭��r�"�f�{�OA���ޗzi,9�[�V���p������[G�UHY�`�͢�*�+4ϖUU�W�j8.����+Y���v_tD"��Et�7�_��*%"(�hQ��53@O!�n<�$�;WYh��	_�\��f�&�֗rh�0
�z���%H�b���M�����`t���O��/�w|@�͝��+��`��'�����:�j&"�8�ݨG��Q��Q�*�J����a'(��x���@�@��<W��U�C��ldo(�NNt��jv6H�	�8�	�*��� �;���j�l���p�츢��"�nY" ?R��킕�>�c�`���
y4X�f��g7�E������Y~2�ap4��2�h���Q����t�!�DSlI��Yp\���cÄ��ItB�p8A�N*\�����i%>�K ���/(=��O����]�ӣyb��
?�X���t�תp�V+����x7�e��dU����Z�uZQ:v�a�r�j�R�c���h�"?�������r�2F�۟�1�_&��q�
��W��gu$���~]خH�@r�M'���!��'Q�f�gN��/H�����
�fc�Bpu���N��&9��L��v�͠i���䆂kw��?Eױf���}�<��kbg��1AĠ@dR�ӥ.PY�'e/20*�Q���7X����k�ED�<���6(!CY�n��)�nz|r�c7Ϭ��A�0��$�1E�}a26nfo;�ڟ�S�э��W�(��O0FB<��I�eu��p����]��<�BC��H�\�4Ò���p�*��ߢo�M�f�"��Zf?8�{:��#���Tk�7��>:�%��D�p��l4���G��@XX��N���џj�5���ׯ2��7(�o �6��s�ţ躄߮/驤�@��j�]a]eu+\X��ܦ�)��)����;΄ ��Z� �d�=��<�H��OgFe�(,!��Z�
��R��Y֬DοOG�)��q"��#D'�|���언?�	�j�OZ�p�G.��%&æӔ��㘛şi{��Оh��L%�jIi5TE�b ��=��6����6���o�f����wI�����>COl-�Ԧ��E|�f�eJkTά�e�G������z�������+M��l3']���#�S������b���@��d�eW�����[���]�7�49�0���ؾ������<(�O����Ih���dG@�ſ�l���ɧs,��HKRI�+�U�1������=��f��7���m��ؽ޴LA"��^���5�/��>�S���3�%�����Rkڡ�J`�̂�������&�w�#70!�@̧#�5�^����I��"B�@^oD��64#�uꅉ�n���E�n/�{`22��sG�G=i�����;�˳��2�l���*�]�ܺ���a�ޚ��2*���3�F.�S�E�cJ�%�Xс(��-!�?�ߑ �h����s��lM����'b���*�)�G}Zy������:yѳ2N8p���1M�9*�:���F;�Ƹ3
iaY���gA6��f�N�oIC�I��G�v��]���P��X�&��;pM�:��5i��}�)~��>�t�	*gc��g�}����v	�%�d�/�0�����f�S���+p�!7�hJ<CL��%cx%G�J}ۃc�n��7��7E���w���8�wo�9�=�O)6�F��B�6��FzK����|Y�&��8�����6�x��am��8�Ù���2���:2��x�Ү#,��B�����Rg'~+7����MS
�U�}<[�t��]9�ƺY��I2��Y��A�B����N�F9@�fS�6�#ME���)���|���`�C��Z���5��cXE2~�쾩�w�k�-!3&f߅?��@|O�GW��m��~@|4^�Y�뚚�yf��xU. f�N(� #�/8pEY�?#bsU
�Y< ��Y��m9��0�1l|���2sT2�.doD�!� =�R����`� ��5��A	p1�J�W�M������B��ԩ�U�a�	��u�x�ũB�9=��Ǘ��(�L�?̸P%���⡶2q$u�/ ~�V=_�0��.�u���}^>m�^1�0����k�v���6����lJn1�%��6"�y�l~�-<�9����3�����쵞'��Լ<�O*g�D�����$�'��٣ ��zTr2. +�%����9�K�I�q��Ӧ.&�B�@���^�Z�����(jJ<]-���zb����r�.Z!3c ɤ��T!X*i���j�*)"*	�r�E�6w�C�0���y?���W57��J7������ӇM}���CՆk��W�a�H��B��Mw�AON �e�L�Sܤ@�6MČi��`Fc��L"E�	�L��^4�.��}�s�z<lF{���Q!���Nebq���+��e�^;� L�~�N['e:o������|)� !��]����m�"06���U�!����F�;���TH��k�%g#���i6YS��~������-X�T_x���@fp٫���6�?������lN�ћ3t��0� 2�4nQ�C�I��2!ݪ�%��m���i�nS��U�
1F�އ[U��(�1��#Ϸ2�� ��]Dm�>��-R깬�e��������N%Yw?�"��۫��F
�q��O�V�&�TM���BRuzb���.�\�[v{��xl��7�'p$
�	�S�2��@7�<lN�:CHg���=*�����/9W2p��|�&3���r~�q�+p��M�4�$�l��d����yAى�����l���村��V�	2ivY^�/��(���#�iA��������qCj��7���K��,����aJ�&���k1�X��Vv!���u�j�f�IL]7���q�5?m�hNf+���q4��_{���L �CA�O�ilW]|N�h��´1��9�J��}K�p�7���`M�Kp�U�\��{Hə1�)S�բ���� 1Z��L��K��s�u� ��⃝�)�! ��D�Ai�L�����W<9������ЬNE��zT�]�Nյn�3���w
'�������,q@�1J��Kn"gw����y�4���ι9�E��(���a��4���q&Dt�>�B��0ia�*?I�P�
��u�w]�k�&P˴r)��|�66�X~,��{Ǻz��N�}.i���*5��kN���p��*���G)��������I�T�\����PnIp�p���~~k�i�[�<oH����*O�%�	��67���	���L"�!�I���TԴk��+~�X[�T��χu7�VlKf��������$�co�F?Z��j&�x�. ��F��s�$�u�P�9G��]��[�il|���^�L��~9x�ȃ���xW�鈔8$����6��m$�:�j�!���S����a�.>�Pي�D�iϰ�po���rNZ�� �t�"UNRM��v�@|Fe��|���דة'�.O�����HA�`���>-T�ǹSsKQŪ;������%�;���&:/��x��e8�����f����.+3ݵz�I8�n���:%M[:����e��\b:,���[���S�Z��������4r΍RDJ�er��x�O�l�~R��X�.�4L,J���}��x_�w���n<�5#ߗ���%�H�.'��E�=���e�Acu���CY������������Lb\q��tN���k���]��E�����ӶV��	�E�gmO�S.Q^�B	>���4�{��!�#����"u���T�g����1��V�Q<ڬpR�����=C KI��i)kF�1f�N�e[%�d<�k�����q��:��X0��$���uB�^�c�L�G�E�>t�M;|�n��p -D�7�����������Z���g:mF�6&X-X��n��vI�O���U���L'�s@�o�5wO�-btt�4�.��_Aj� !�x�!z4�N	�M�f�|��2XΆ�N� QU�}Ť�BU�0���ɿA,�N�rd��״'mLV��	���s�dO��?�鈌<�oS��xC���U�r�$D� �߇��;�y�r�A���Ñ"Pq�1���t����1��;Tߺ%*`:�"	��a'��<#��ͦ5�jv�b�ڋ��g�z�B��#���`TMpQ�+�Q2/�A;s�*e)*�#R06j�*��Q^�\j�`z��	��v@$��u�8�Sێ��Χ���ni�6tke)g�P*L��K�<���:(�(�zo��-lNs��0~p��.���e%�x����Fw��yW("�%S!���`��Bщ�_YW�Iv����Qw��b�v���m,�F����|��%��,`p�$�Q���uO��t&0�&F��:�x�*K��J"����V.����E��g��u^Y6t��`&a��7FT��G��V+@#����Z=���M�NV8�3�6~t&��~v|م��V�	�z� ��'T����M_��B;��eY�r���z�Բ(����d��)p�]���y��+m����J@���9�S��5�k�4��X\��_tފ�+'��̦�tF�y����f��6���A:���læhԊjd��*
$1eh��՝�ΪP�#�s��Ϧk:s�p�n�h��2�ټ�޸gAH|��l�l��_�����L��<,��
ǝO_�iFe�0=������E�I2��
ۊ����|��Ly�T�](���п�v�o±�Q5�%7��?�؍�f��FX n�f��p3g�?��b��T�:�M7��i���Z����g���Ñ�>�(�_���9ݯ�x����o�]�-kR����~j���ӟ�P8�n�d;�}�:I>�{]����U�'�����O!��"�p��N�ă_�ebS\7�I���7��ѽ�g+I,ʎ��Ν�+�;�F��J�'O�M娱��U�	f��L�w��z���5�M�f#��� ���d��EdO��*:!3�2���B= Ĕbr�\�U�"��bj�̊�J��`d�n����yBd�M̧���..��;�n�̅�,� Cj��il%V<N�iz������$(��j�O�1�6�E`�%`@C��N�+'��v��m�����ľ�.�,����bR�v�a����/8��] }�w��{U.��)[��ETW���)��[xC0���r?a��B���:������`��}_�}��m���G{�pl�l�Yu��qs� ﵊`�-6�\N"g�~�_+�tL$"�r�6��8���{A `�m��@�B����A]��/i5��ӌ2��ɬ+ �I��V'�gCb�Fǉ��F�f�d?g���f���
EPLuB�1��B���Z�xמ�+[�?�&����JR	Ǜ�qo��#G��tV�*ڼ����{�'��%���oX�U���y�%fvD��/��7�F{�T؍0w
��	�(�T=f���<$BԺ9��C�>hOo ��$�Q���F�̲����k�蝳����%���ӹ*=�C��j������ALa���"�Z +8�>7�m#����YJW gDr%�d��81�/;���G��]��v��f�i�?�JI���������3�� �RZ�3W���#��,uD�aU��c�mK�&��o�i~Ս�S�M��[^�\ޣ�ı[��J}�h�S���؞�[p�̵3*s�c5��>3+�6q�翣�l'��P�h��3pS�9q{oVx���b)���V�=�<+�q�O���P��Q7��5'2�)����8Zut# ������+\5v��ポ������	�в55J0�@��U����y��B�Y��	~��*x�T�?�b��#�}���HD&��X�R��b��Iq��*R��ފ��Gr��`A�:^����L����,~+,��k�ˑ)����ݝ����:�kk����I��د�ꓸ��9˩����4�`��*G������H�d3���{�þ��TJ���8�$¸ӣA��w9��!�~��FI���6��Mi؈ݠ�X g)#��r2��R����|p>^4�K>+Zz�A�����n��"�0!w���p���	�/�*K���2��*�C�|��2S�+2G�C\����m*{���ʓ�������6h4-<����ǠҒ+v>>�b��>g�{��H��'Z��PJ�	���^���rbv�xG�}������imG�Vm�H�f2���O"<p|���Ƭ��}#�)x_�#������*0�ML��o��2c���W��v��R���xW��l8nĄ�ɯ�H�[���g��؜z��  ���B{0ժ���c���n�R�B.p>�m��L�ͥ�僢EE�a���׊�KK��>v���4/��G7u Y���/"�_�v��e}=��0�2A:��&x+�%{����pV`q�X >�F�T�͕�kEH�������k���ٷ�,��44�؋��\�߇�^���H�I�!�\S�0�di$�����AWͺGf�L޽�U������'�א�'�����c���"�~GnA�?C �?�c�rmI)�f�x�t����C^+�k�<syI�<��g"��&��7616�� d�Ֆis[�Ib���w��&e0�a��H��~���>"ཁ����S3�kw{� �kj�Oa�F,�-�0Q���Q�6�Sb�P�}xgQm]B�����ʓ����S�
�|��&2����2�]�H��u$�+T��.Y�¿��~�n^��?Ag�d��|é+?;��r��r^%m�YN�忲8n���N ��V��xv�o�2�z%������lM�e�V�&�&��c�UCы�T�C�?�є|�蘇���p��>aO$H'h���(A��FE�6p�UeM�d�|���������c��0�|�Q���Kr�Np����3hc��R\!�4ٙC�JNN�຋q!�6�LU|+���O��zХt���h�n <�0�I�!���q`#쟄���m�9g�Jw�XH���؁�t�$��0������{@tOڞ*�#e��8,T6b���h�l�V�pvx�QV�F��~>t��1r�H^e=>���ɲ�^�7��z����!���mJ?	5�3�#m�"6?���������?���31������������g��wl=�H��F�(�]oF��"�kҪL���4��T���&T]6a��,�'����D�$O�%SĖ9�:G����q���^sEe -�g���@���K���+��A��Jx�tR����b2���	�7Di�Nr��Sn�ڜqh���UfL��fP"
������F&�Iߊi\�����I������~W���{�K�N�|��s$��D\��xp� �λ E�ݱ���WQ�o_(����� xnz���1���֍Qt���dÔ�m��|�̑��9�I�1'�l���E��P0��l-Sֵ�����%���W5CCm4Q�րG�s�%��w��+mjeץF��w
_-A�h�U�ؕ�>����-�
I��/mzz���K0�h�N�����������ND������KP�Q�(t7o�pV��SR�t��>���s=_"Go;f A �ᢞ)�t�
��	���;�Kc9,@J�S�"41�:��Hz�����~���Px>/������t\v�K�`�����u6WqZ�&�檗���҃����?���U��;�!,�:p�M���WF��sT��0�.��}�"#�	�ђ�E*&�+��Fg���hq�\0��]}3乽����N-ԍ�� ���ӷ�����R6�M.,,�s	BU(	���e;��U��� al�Bx�Y%b&6��o�(�7E�[���If`A .|��(�)Α�'X��؎k��Y�u��JKkN�fV)±���Tl���X}��MZ��}�.�m�r�q�N�9��?�f�h��8�a�o*�Z�� 	��낚�B!��u�����]�/tcw�Z2�g�J����KƂ�RnU���6�
�뗑`J���U�zb�=@x8 +T�ao*l�^p�T�E�*�Ug�ejE�x��
y&��8i�U�򖻉���i�EQ�Zh�nz�]�cVBdAk]��,6T�Ssㅡ�b�k 0)zaRB�Y]{��v^U������=�*C�P��x	�i�}��<0������'K�s"=�o��X�m
ƭ�zDK�����W�@n+�lC��A��c�77Z��H��So�?7���_����%�q��l�}MAF��^���wl���,��)=(�Q�����~�"���b��Q)��s��Δ��m�ð���ٷ���������j��0b�m�|+-)��:��ˋ=L�� 57ִ��Y��0ڱ����w���㽀�X�y�I3"�(Q�^m��+A��,��R�����gD���bښ����O�R�a!'���+�֩�d�� ��Da���W�������~�;�3�׫��N���A��������IOy �e8?�����+����㖏��n�K| 4s���/f��^���Zss0c*-3%��m�ߵ��!E��/�vk%�`_xٿWg!�o �U�Y�t�ce���Օ`�t�|:S�5����b|��^O��7�Ι��`W�Z	Ψ�.|���+��P���j{a��!��L:n���xȦ�_�iV�З��PтA��nq���_j<+,�D� 1*���qә�9m�e���]����u�6����?M�Q~�m�j(���8�`Ds%��9 9�୴R�+X%h?�b�wEG�J�)����_7޷�#1B�t��}�������x�/$��D Ðx��U���		Y{{ �=�u7�l�l�l��2Mo�?e��j������9]���a(�iav�֩��"�C�r�Gd�p����������G����I4���n����t:�V<׬����k s��Ұ�����ԗ�2���x�Eܵ���[� .ws��;�Iw�s�"����������j'�.����Ey��y�F,�O0��F�щ�>������^�C��[�����tb����Y���X�"�F�1.2]C2��C:��9S?CzmЛ�R)u����Ae�Qfq��l�i>�p�4����RT�g����Ndl|e���7�_8c���Rd���!}hC~�����{����a|�R���B�Q4�ߌ�w>�:K�<�l��E ���[8��x����cb5����I�!�rv��c "����7�:���^Vh�S��޽y�r���[D��]H =Ш-�4a���DL���Ds<>��ݍ�hE��ӎ���=����4�EQP�h%����<��ݑ���VVqג�����S�~�#���?b�	�����^��n6E���<���w�>)y ���Ϝ��B����`��x'�,2�a�H�L�B�����E��UӚ�܈j����ߞ��=��z�\��_ŨL��ct�N���4����S�w��e)	��ʽW���O&Oҙ�~�nQ��5�`,v���3IR�?O��_��6�^4yH�.^n����?�8W|��[)�=��������f)�g��(�2�O+�����`4	����>���$�;��v����æh��& �%�(��A�4����4���\od��]%Nn�>X�>��b�"�u@��Ζ�qM��E�p���e@Ղ�z�d���k#��&A��5��^U�f�����}�H+-��$@ѹM��
��� ?Zj�c�^�Db�g��l����3��-]~Ig��|o2�R��o�,�'���r��Y|Y��AJP��:�b��m9 O_����ź<����T�[�i�+�85����`FOp2d������d��u�ͦo�v���p���B��V�!78�V�&+$�6�H�ƭn�za�*�I����⿼�A�W$w������ȅ^�g��<u��G��m��-��3p٢(��գ2L�Y�6��,0P�]s�,���U�,���������dJ�$Nb/4My!d0W�!�6�x��lwUuZ,��\��?���� ��^Cǚ���C;��k,Fo1���b�\�p�mE��S�#41��@$ޝ<n�ˁ���I_뫻q�}�EA(��`�9�4�K^�aB��?�u �5YE��m�j-Y,��G/���`�n�`��S.����]pF`�#��/ �����y�"�ݠaS��u���"Pe��'�'���Nz&��c(�\["��M�׃����za7�9+[z�g7���6�ƭc�]ni�xBhb��nT3�����ꈞM�O�Ì������I��s�]L�R��G�$���y0Uy����=�`e�+��
z�>����x8N�m`cI�(/y;�a-�Cۣ�\�`M��� 
m�;(10�;a�/���?��(16v}ʶ��/T�N}'^�H��|��s��s��)\���ݐ]I�{F�����d�Aa~:cV��k�&��N��W�����E� U��D�N�<�/,B�j�6�(��>���k��lU���G��ؿ���n<�JQ�I�dp����H�\38�&�8��t�R�~��&�I�Df���d�B����?h�%���<ʈ_Zj%i�8��t-�	�iP�?�NYw}�pY�3�r%U��L?�^{��NU���d �n����8���O.�t��[; m��^U���8��N�����m�|E?��*&�>�\������([᪾��M'��ї���dD3ʐο�vŧ��@�0�`d���ڌ��Jh􂥭7��)�z��E�Yz:z\i)��/�gM6�tP#6���D-����͗���R�Rv�+O�E�@@��NK�Ey��XpB�	�|"�����SoK�]Oz��e�9�(��N�U�U�&���1�{��JmYr+���+�AF[+\��\�T���k�m�F�N�ce ���R��;�kl�AC�����ش�����9̕p�M�ٙ�����$��I�14>͍��C�h�Z��/�G(�%�{���P)u�]e�zu��(k�$e=�V@�63̲��~��^������H'�{ ��?Ȯ�����zٻ���h�G��_�2�շ��9�I0�⤦�e�*�´E5U��䠋����]�'�ӠF?x�h�S��0=�<� ��H���S䎨�Ĳ3��%<a��=���X� �D�cS���R?��N�;ֶ�gl�b:9�Q�q�y��)���ty)���J�<�-U2�oí5x����.yJ
!�j�X���,7�'����@��G�����_�X� c��:tk�`vo�mT�͗��zR98�&�v�3^P����x`���� 5NZ�C�t̂؄�>�
&����t�{}Rs|0A�+��YCfvI��T�Y� ����x�������\��Y���� 
��c(�4�|MP0UG��|�2n�f��U�ޝ�11�m_�����U�����Z�[1��bC%H&ޓ`���@ᩎ� ��羢BU޶�)�iQf\�x�Oz�ݻcݤ~,��7����@	(�|���)��D������4����.%���L�����I�1x��Q�p�'IB�_v����T}t�.��G�"����c�e�V�	#��T0�J*(�cJk���L��T�:rwz�~꠰�Q�wE����l@�LQ�9�vE+
�Щ���=�>�u���%l�����`O��úm��d:z��lC�f��on��!�7��̟�t�'�`��n���[��g����7	>�I��ZR�~�.��ճ���f��W��m��m�-R^$�2W��	0 L"ծ"j`#��[��I�Y!���k^ؒ�p�k��]�dLd$ ٣���~�d�@�Ip&���9�I{�S�kX%v�L5Y�4��|L8�/�Ϡ�����~c?nO�+�R�,�Y�l-�<]�M�+m�����\t'|�I�f���ݒ�W���+�)���t��|�w�-�b��Xo�ώ9Yg�����Zk�!��e˩���8���K` x�%�e�/� ��B�_7p��� G��1B�;S��U񅑰 O< ˷G<J*ܓ���B�(	�k�JB*ܭ
�B�D�9B��}� ����cT�)��5v�W�W?�n�0ņm#Π�w���ս/|�ѱ6�H��[�׶�:Gm
Rb��I�X���γ�x�\��F(�|Ꜯ9��2����Y���o��?����>N�R�,� ����47�#|7K���KX�G?��{��o�{%5^��*�X�����a	,�؀w3l���qK��P�IR�P�}5C��f_
��*,��W�7 ���-n�czq�?��`��̔&�cc�/Xj*��W�*M�<���p��j���U���}]����/a�,Gq��诽�5�4��q݋A�����u�3O�")#�^�Q&��¡ ���F��U��gk�8�͆�p;�Q���YjM8��e,ʸTR[_�G���d�&u�9�F�J�{�(m!C)�6��F�E�
 [��Ud���"����/U�+�`r��B�y�8.�A:�«=�l��+}1>d���^ϚZ	͢���p	[�Ў�=>���m�#s����P��.�]�9��Ћ�����;c޽^d���ׯ4��a�#@E��Z �Nu�����B�/��j6�8u((HV�l�K`��vD��ЭD�"��'���3����D��Wծ]5�}�O(ۿ�\x�\q3��p�^��B� ����9��@�ܴ�{Hy��-�H�b�dN�G��+̯�ɓ<������/an�%��Q���u�'��7wC�{�!�ë��?ڑ�A����1����3�������O�L�	��OC)_��Cixݍ�@i8�	��Kw't����Ce��p�������Y%�yY�x!4�Ɋ��lվæx���)���z�OQ�"�����g\h��>s�0��4��/���7�+��h`�t���TXS�>��]���KLV�u�e-�q�  Ufs:�臫��\��D���1��J�@j��+=hK���6�S�-�>.�s'���*���k|AZ@��Y:��QR`����a�CQ���(��GT�F��t�>z�t�u�Kp�^w�
Р֢�#H-�����I��5��z��gR�?��[f����X�!+��$19�y�]�35�����{�xt�/�U�z�'O)��K��sC�<{5"d��<Z���oSW�?R�L>��j*S�'sQU�b��c�yA�s�p��h��.�&�p������D0$Z�K��n;- �9��3C�7��X��㠮����.��M�u܄l;4[�G�F���f�U}�8��+�^�osV��qH�b�-ڇ]�%KٞE����Ф���ȵ�kskźT���ORV�k r��֋�.�2DŘ��Z~��FB�.�<��L��2���4�=iq���ע�v����g;�ٱi�Kkx�9�e�PF��;���	�|�x�l�5$��r̶��QX���:T���Cፎj�&�����*"��'��ف��n�� ���q�~ ˼C�+��'8��|�5sYR�d�g2�t�qzل��x5���Wl�(['�&�i�s.�ZCUe�����㍿���OE���f����b�,��T�N�5�͚q��F0I��8�8�	? 9$]��y�����ڱVe�X����a?8�g`��Jz�b�d6V^':t\d]xƚ.u ��
:�d�Q頡�o����EG��u^���Q&�(�h;1P�H&)�XȀ�^�����h����=���vK����!=7�$
�^|ѳ�b��ܱ* �8����]��6��b@��'Ǌ�U�4�����e2p�
�v^��0̓�}H	�KS�蹂XHYU�w��f�O�vR�Վ�R��g��iLhR�9�_�ة��A`ٕxzYt��"!:�],/Т]���T,�w�`� Ȍ� ��ۮe:Kۘ�鐨�C`!��1��,�a�M@i�4�xC�1
����=�W��N�����~Y�R����1ù,lc��6"��3�� [�	��Hu����C�{�G��@+��UI����~��n��0J����D��:p���d������FJ�t�A�+��	"�*Pc=��*]���=�f�N	��m�o�eߚ7Ã,�ș)a�i�A����vs���ًmݨ~����� ��Ӻ6�"�k����@�%���6�鰰���2$�U~����_��.E4vB8\3�V����nc�e�J�[fp5@�骲�K��tz�)�.	5=��\;�v^���<��v^7��T�&�s��H=��R�R9r�L�L���`�B���M�W#��O���B~�u%I�����<\�S����,���F�xS�^7�v�~F�ud+_bX�A���髟.cn�s�#�L����S���Yi��_�a�½X\�gs	���IC���/+�5R�ٖ��o�`��Hl���t�.e��<�(5p�EF�0�O���|ci6=�wU�!�g*&���WG� ���X��� /{'ڀ���@��s�e�H
�P�fM�hН'NXR`�NϮ�0������j��SmD)�c� ��'l�O�qQ�b�mADT�y����k���C��0A��$��8�^�z�>ù���
k�R"��Jcs�L=&��>{&X�����O)kfz��`%F�P�;2�f�޻�U�^����$�%a$u�����%���bgW�� ����]��:P�!\��j�zk�4���L`���/e@�RC�;'C�[czY1d�"���7i�w�l�f���}qt}��L��{`Wb�c ����!�Z8���th��M�(3�;C_2FtI�$Iۉ�9��Bd��2��`����5Hм$��BZ��mESF�0����s�d-ѥט>A'Ȼ(���J�53����V17���;���3J/�Y�I~��Dl��K��-V�"2�+%Y�>������B{��"�w����1��xe��ݴdb��3���a�7���޸�Gxt�jI�%����;��c�i'�)X�Kɐ����5�1{
k�#<�ζ���n�>��*%by�$:yjy�r/�H�&��YG��f�u �g�6A�skZ�_����6]�򢡏CGk]޻ܻozAR���2)\)ѡU���CNF,�k�'�%��f;�����BpW7�[�~ɕ��K�}�Ƥ`�0��%_~Dh}.l"�\����o�m�ld4o�����(�T]�zAn�ME�YܑW}?�����y�����S��hPD�˽<�3K���s]u)H�Z��%���ӳ�@���>���Q�bHЇ�j5k�`2�V�p���s�4��V��W�]&.-���N�??��g��Su�m(ʒ��r��YZ/��SG�V.f�8ʶe_[��Qc�a}��ϻ�$+���iօoF����i�V����K��A8R/�!���ؔNؗ�@7�2�-�Z�v�P ?rEj{������X�kj =�h�:�&3�����&y�0��i��=��!p8� H	��O&(�����܅��K���'�0���$Vmr���a���K�=w��9��/"��x7�qpYBy���>x�!�����f�HXz�F��)���^�@/ԡ�	��>�, �w�� fD���1\u[,�`wR��\~"��EX�%H�k3%:�R��R�>�>W�?Õ��Ȣ���^D��(�ud� ��R�b��]��n"u^���}B�t{���^ d}-��[Ȁ`��DBE��&��@��(�� Fă�	�$�
� 5���Y�iE˼k*FѩUۋ������l��Cd5m}[��� ���q�����d�*h��`�,;��f0l,��z&�w�*���@�zuf/�	�2�|��:&F�l�� �H̪���$8u�/�U�)R��#oؗ�w�0w^ 4��4�E�O۬s����m�ʿB��¡2$o�����ޱpA7�E����|�(�q.�����k�h�]��9�4��L? ���B���W.���D�/���1ův �Z+v��ã]��ـ_L���2�w�&��/v?y��x�a���1�;0��U��VL�y��0b��f7ʘ���ip���L�����-�,���$,�D��:����z,�P���cx�Ϝ�f_����asC�����2��C6�u���;�+��õQ�(����<
�m��M��M�8TGW{���U�՞ILqSh�Y84N�@̰��c3`蠌I�����ʚ�Q��c���qq�[�@�P�e {�$�s�Ȝ�v�Iz��Dh�&���f���h�Aʝ*ù���+�l��l�R���\z��F��ǰL�����}���Se{�r8����TJ��̪&��%2�� i]�¡8�������������/X3�zE�0��;'F6W���TkI�YE ��9o�/:�Wr�Yf2'���Gk�������Eٖ�!�G)|����������'�~�HC����^�Y�ow%��d�gm���ޗ��gd���Z�imr�4D�%~���]�'��j�� ��-�R��8ĳ��d�iI�@[>@��Թˢ�v��������FT9�^�v�|9OsA���eL�ȉ��.EO����d�*(9˿H0kD�#�����G���Ռ��Jp��Zi��� � ���4��b����$3��Z� ����>�׆�h���O3N�9��]g�p��QT������f&qb���?pԚ����/�v�/O���
��&xYe	(�e�;�e0�S"�{ýsm��{�^C�ˍ`�]e��*�ˑR�� .xë��@�["'�3�>�N��8�I�<�y��|6K���p3[�K�˼�6�g�U\����,��֙��9`⮆�p�O�r�W$�q½ˎal�1���1W��Y�n��~��I�a1�	�-K�5CS��2*��T�(|���o�`TS7-L�R��~cY�k�:��L���a��[��5�m�Y��X�fXm�]AE=��_��|H�Div�L�Jc��4]�ЁA�S���'$]��ӆ�o�i����t3���Q%G��T߲��o'#�����9"�1h�٣�83�W�'��(�4���55đ���i�����C���ܬ�[�^��Kq�N>�{���80ʿ䐭14��EE#��©OLQ�3q��`P�@W�.w1�
.�Ή�����wo���7~��쥋����A��&��L0RV�8J���6���C��r�	]lS�6�k�vk��7�c����;t���>�E�����j�]�`'\)����RخV�K��Z��i�'��|�ɳ�W��7l��,�0	dh�<�T��F<����
�;��2i��!�L�Ag�'���3�!�D���Q֢LMN��p��|�x򻍡���>C��D��8���g>�p�%�"Mq��(䤂_:�(_���P���q�@W���-��c�	��r���V}�y������K�4RO�jت��Pg��.K!�}�P����:xax;G詫���&f�F!U3���)��y1�t%cR�;��4J5�i�lG͇_5��֞�D]8��	ǅ6n��cI4�?���3_��YK,��r�6���PP�0��u�<#��ƶO�m�k&RM��{��ov69��9��i���З�L1HR�ʞ#����g]�N�t�J��x03���TY����D����3YN2L������AG�?�7
GV:�pB���[�b�������s�ԫHy�<�����ޔ�;|��4֨(��\��6|�#�3v8�H'�k�n�E�@Z�D��4f\Z�i�B��yhEX�.h��j�����Ѧ�ϓ�+!t�k-M��D�|^ z�I����Dܛ�ի������
;�O�(~����h��3`�
��\;�Ρ����^�~g����y�ȴ�]��G���5m>���&P50{O��p��5�b$G��5�`m�0��������e�"\>��m3�b���A�F��M��F�V|�[�ƴ�Բ[��UX WS�#�h�Y���dni� �3����&���R�N��L��e.-P�U�;�)�V��a��ΐB.UwRmQ�i�]�
�c���Rek���Ѕ;�Im��sɍw�!Q�\�L&^�+���fm�
#�8}�
1,��9�-��|�0��7���j_��(k����:S�`(������z�a!�, ��7W�J�i��M9�l��9x��G�%jf��`v������$Vw*��O�J���@K�I���B���Q{�8��n6O�g�¤j����s_����yFS��P��i��"w�/��'D'Z1a�]� UQBJ��ڴ�I�$�C,�0v��|�rҖ/3]9�v���~�5@�D��[S�p]A�y "�8��+E=�s�.p��I+&Mry9B�p?��T{�5���[ܒD�'�8މߒ�^#�i��/�;ښ��QW�V1ϑ���\��ږ��w��#Saȿ��b2	1}����0Sӌq%I�u�s.5�B�WL{��ƙ�
��d:E�Z�E��.㋮��$hO��,d��!�%�C�O�e��תiX���+e��\V4K�'W��9��W�a�h����Fa5;���L#㭖�5�pHC�Q^�ݟ8�xד�	�� 3˘�y"������d��%[�E/4���ޢۈZe��`����T�ܐf�\��/��{�ou�ѝ$�#�C���4]��Ŕ���5Y�3M	�\ˎ���4�~�ךZq�hz�(���O'�awO�e����<>~��1H�'8l�B�H�G����!$�i�!�0�'���~R���� �d����qOC����a�6�|�	} t�(��^f��%m�	�δ���A�>Owl�s��4ϧ�λ�d�b�d�����|�l��rS8`Տ=Ȟ$I�^$\�����`*��J��3�=���l@��s� �:[)5��G�IC(���8#��(���bb�s�EϷ��݁��/���t}�,�Y�Z�V��Fi�R��`��F��lĚor}4��*�,\7_�C��:���3�z;�r��r�v4��%�7��������S�<=��p����d}�� b>���*E;�L���;u��ey�E�l���L� �Tmj���E ����j��hה�m�9�z���[�$�{w� �ڪ�J~���S���Ns�Ќ��-EHs�N�^��X�n��u�@���3H�Nt$�5�}ޱ�,�L��(���p2�\��3��RR�J��7�_��'�H��������1љ	 ����;�1��;�]���d���0Qs�̲��Ҷ�_*|T>k�'��K�RJ@���4�Q����,�k�fՍ����)Z�kF���;�c��c�$�Ό�Kp+&=�ާ���$�_
�=�ߨ�a��H�C�J�Y����1�3�����RxlO��@f]��M��v\N�^����Y�82�*�+u��1h�������+�dkR/�<ݎ6����������4������Z�a;vB}�]'7��;��T�n%h�߽ٵ7Zx^U�g��(�n�M!�Bؚm)�9�)�ӿ/�x[��aڶG=ޫTX�r�>mFH�{�W�{��ۂ}�x'HK��2�p���t����=��鴲`z#ý�=�;Ve�07�!ʱ�O��]������`��>�pcO%����v��o�$,mݷ�g��+�X��x���a���W�_�ۘ�\(�?����}!�	��`ֺ�[��iRy������?۠泦�/����%�_����o�N�s��A�*j�&�p��Z���*��A�a*��T�u�Q9�+�&�^�2��	1
��&V5!+��2Fv#�V*0r���yW�3�ϰ�7����L�l8,�kB�C��ktu�*�^X�_+��6T��}tA+:�l��F�n����r�ܤ��i5?�%n$k���b��ޕ<ꯑ�I��ڴ��
��㱊}��Y��%�}@��J�</[�r�����LB�u���훵 �C� ��� �STF��Wn$�_x�ɲ̷�&A �b�D0���JFv�,�S�6P#/�z�o7 �oÀQXB6�]�Ӛ�?�4�� M���N�;]��t�u��l�M����,:���"T�FB78���`�`sh��S7��K�L�����TH����\�Y�I�(�*R��nԅ��RO�����2�C�Oύ�F�)zA^�+:�:�ޣ��bҧ���&�d{��9�^u;%
E��%
K���P���>�ڒu���!�x7ж67�C����`�2Ё'~!9�������'��8V�t̍�M�?�F1�@\?-9>��BZbo�Q�a?���I�ĕ��R�A�	��)\,;��)�Yy��� �6��5\u�S:c��/�٫�0�[c�Bf¶�U	�����p1/��w����_Vr3>h��7O	Ủ'��}J��V�A�TtSY$�I�X���Ƴu��6a~�'ü�W�/����Y�c($du	ˤ�����5�qgG��',�wp/��|9-~��|�Ð�J�d:���U������ۃA�?�q�fe�����ԅ ���p����92�Q��~ÈD#��!e6��UT�j��<��$[��4�(�`���W���7�\�����5�*2�
Y�Z_�P���}0,#@��i"��T����jJڽ#��`k�oB3Ky㘠���	�+NP��;�0YQ�8�݃%vT����gs���̛�s��{*3��U�|�z���ɋ���'�('��|��\�~ q��BV�m��Zq``�Vm
����m�a�>� ǝ�پw�?�0k6���pzp-@b^�r�/��|Ș��mX@BZ� �r4�ÙA�f���P"��oT��͋�����G�}?X�X�}�֖����d �lY�#��s���*DKI�0�L ���uKz�iJD�`ki�Yq�f\Pz�:��Kل�N!�KLźV���_M�F�c���8;k�V�A졫���gSL{��_2$
�)���	In�!��O�<����'0�`���7ʎ<���]pO�����L�-Z��`R�7u�[�=@ ��{u$ �A�Ԍ�5a�j~cCI�|�Ť����xғ���x�˘Ѩ�'�P���O�3�;b��B�^� ��"��C��}M�c�c���e�ӷV�%"�h�b�s�]�=^+���ۉ�g��'F�9���Ô���cb_���̉�%����$�j����d�%c$�F)sE�^��Y��zO�܂Cne�j�Z;aw����U< ��l��2�BT��S?q(�F��5��n�o+�3��J�r��,*� 4�E���V����ǳ"<ؗ��$�����54W�U�:��,ˤ�)xhbCc�?Kj%������[���/���X-�����|4��)����a����ĺ���F�,���>�l���{KDP��vM��i���a�,��(�^ܿ����Nau�x���Z8�T�/�5�T�����滛��w�z���'��pB'D!u�B�S��Hm�=��):!����
�����M�.^���H��,S���T�W7P�������	TR��P!�X<�>�q�%�G�1.*��'oŶ������)+�y\�ųJb����S��񄅥콓�?>�t���Az[2���̣�=s��5�͛��tݰz�|����:;]
`��Zu�jKdi<�1�/��"��L����d7� I���� 3e�¬�����з$��j.,L����i�@�[U��+�o�CI�S���6�H;''���*D�����3�̐��b��8��jv�Qa�ь�; �cS�O��Tj��Ye�c�>ZhAc�o���1�a���3q��>*5�����T-g�U�Mp�i������dH���X�+8��Xf!*@O,l���J�yi�����V;�����K/�PE>�j�f�zZ\�8��M%(�f�����4����Z�H��`����ة� �ӁS�7�C7����|��B�h��&�4H�(�6vk:_⩺|�ot.��W6�1Of�74��T>dx�7�=O���7ث��>	p�nTU���CQT���?`�VOAnڏFC�$�q>q	� �JJ��Jdں�c0�Yb	"y�{��:}�&�xr��7���%��hk�Mɪł�B8 �F��C��N��_F���;{"�]+UMZ�`��,*rї�
<���Y��w�:F�Bl�]ui�B�B��f��C쪋���s��	�D��>!���	�� �@!�Y�Һ�����z���+��	{T�=��z!i#��{�3eQCa3#[�e�+t��2��֧+��������~�Q#5|���c������ʓ�WݛUk��9>�Jl��Gf�9x��Mw���;�eP��T�2`pzE���y�Qpd�|F HT��Mŭ��֜�{{�u�����?�mԢ���<8�P��!s�TpӪc�	��	�4^�/���G� �P8 �r��2w�"�T����	����[�n�J�V@�G9�}��T��l�K�/q/(L�zz��Jw���O'lp
ng~1�+U;��r%?����
�1)x�_͘���p�l���tW���>vM�^D��}cD�H0��F�:�SMLRcF���=]c\�1������A�	�Z�+�ٙ�n����A���o�� �ku7ݝ��e���=��>����	@�
����H��[��g��' ���
'(�Н-@�T�M�5���$9�d����ّ5m��@W�s�[�&����.E.�n�6��i��w�㭶#��mkD�]�.�
���v���zȴl�SC�{4�=k�7���\�8 7qE9�H��,F@"���q�^�J2�w�aa�T6ͧno� M�xʩ�XX%a<��byvn��G|�cٱ;-����SπBt�S��J�	���Z�CV�`;.w�
��2ݦ"�Kr���*���WN�H�&�8�t����[n'$G/mᢎ-H��^/�Q���"g~�ܐ&d�bWa�=L�x �G��#5ځL���b���7���(bG$��{�Ft���r.�\ǟ�Q��|
<����a;��V)ln/�tD���lϙ�y�R��)D�Y�Q�p�\lv�����t�2�:���a%]��<��S��|��ύ�����f];jb�])�8e��PvY3"�8DUZ��C�ao�,^���<�8ͺ�P*�^�ń�|��)�0��t���O?�M��O����%"��e�r��܎M�L���ݺ�>+�Z��\�k:��ݚ9ߛf.��l�-Չ�&�d��� "������H�!���ܘ�I��/U'�u�V���3}���V�`��x� �%)VS�%қ����L��2mu��'��ͦ�X���}�MW�������u��%��#A����>z2"G�/���Zҭ� �4,6<�]\�~m��N�w��|�L[� g�ı%��R�[;�;�:m��٠an�W䧝��[@��|h�w��R�J7�E7L)N.���{��k�`��e�N�S�x����N��5q�Z�7
&���V��̱���+�XM��3?��۸��"4�'X���Q
��M�>��q�x�r'[��W�^c����.*����熚�� nGДQn�-�|��V��� 8�+Fދ��b=��joɩ(g�S��� a�*��`39{]�e�M�4�AϺ95V	�	�}�N)� �p�6���Ju�N-�5�~.�\
��s2ga�=
�'�;[����>������b�k0R�D۶*�oF�p�p�8���8�~ݍy�9����8�g	���p�<@��̞$]��mE���k��9�>l�a`4����N�����q�y�:�H���挰 �"�'��2��m����0eJ���+P«��*�X�[��.X*此�B�&K*;�p��2w���?�E���VH2�o��_��G��2��E�׊~�f@��vZ-z�G�]+5�D�B��t����3-�}rq��B�r,x��II��-�Zd�/��>�[R�U���w���Ji�%;�yCX+�]�5_vP�ۣ=־�z�����CO�T���4��׽1�6hB�fb܄E�S�WB:�}��P�=�t�.��wP/��4���80�Ŝ�C�����Q��A�^�e�u�Z� Q�޸���N��H����}=J�TE�[�Fƕ�P�L?�LǵB,��ٟȥ\[���e��s|���U7;����0�ޏ���!ĢT`%W��a�4󫔝8�(ȷ2�mXY^�*gY����g���85m�|� q0?Ǚ ����� ��.�CpZ�R,������˙2��w�3�f��bl�SXsk¨�Mw�L�D�H{ɛ�[�8���t�ɴ�$�������>j�q����­2������&A6�DvM�;�Y9�����������b�@��i�����j�8QL�'i��W�s�����V_���Q#+��_k��@e��s���5�1�]XxEBk�s�u$��Ҵx���;�9�NZ(�Vscj� �<el0��,�Q�.@M{P[g~NK]����~�M�Sjq;q���@�=w�4����b���mN��W��]7I@:)ڊ���.$���x���H2ux8/[?׃76#:ൕ$d�?�ҳ���J4C���3�mе��1�P,�`�b]V�����L<�Ӥ�?�A7)�Fn�n4m&�>^��u���_.�k�3(�V�܄��U3|	��اG�K���C�eS7(������o�*b�� �.�P;�jF�*-hj�RTݿ�!)6�8�D"%LFc��	�7��6�`�aj�sS�ۆ������ԷՅ�Ҳ
�}��?��}}N4*�Υ2[�4�ڎ��
8�Q²��ơO�@/Mᬺ��kl���5�F�x���N��E���5� �E�C6ky`��R����`fTHjy���J�p�N�6���$Z���Z5���ls�!�WCH�5��ZsD?����0.�8q'�Q��E���5����%�o���5��cߞI�p�,DJ��j'V+ܯ����/)���7�,`�V�Na���t(�u���E�Ӏ�y�뢆�p���s��	�I;���uݿM�x�#��]��������C[h4$3���bGd�@{Z�/c<R��+X�Y9QC�A�a�F=';�T=C�M��ü�_qX�Wv�9B��^��c���������X$����B�[%k�$��oT��h!�I�ǖ��v�3�Ӧ����q�.�A���G[��l4���og���[D�k�Ђ	-��,̛	��J�9[2)�&�+xw�b�լ��f^%���Qk���)�V�t�g���d�;O����k�F��Es �n7�X�c\�_��D�-�MXKR��u�ihnG�ʋ�{~ �g����e�;6�c2�����H!��vM�'&�ҏk�n;�����Җ5D���(v�.6 kI��������-Ӟܝ&]��{�� ���X�~�P���kЄx��7�}��ѻ�6�1]�9��KDH��*qv�4ݓ��v�P�Vd��`�%]�)�[X��A��^�]� �s���W^]h�W=�U�o
��1�6	Z�k����*��yJ��<MK�eZ6n�.�r&7�w�(��9��lpw��Kv,=��ON#����H�;>T7�3��M	GI?�@�����M�(z.�	8	�j<.(H#����Gw9��h�J��UG�=AkOT�T�RT:+]m\�C�\��N`�.EwX?.:��M�eO��]����c�~`pB87n��7i�ڍ_�Q��m��r`���La�v�V�����d(?�p<)��C�O�'vPfƊY��`�	+������>Q�%(%���赙sQ�-i3�v��"��Uk�+R��}�B��)����3��lܯn�$�n�/��%����dQE�$k�2?���Ez��J'�%���o}��-�76e��C�8�;�K�f��3���kt��r
��mr5�A/6=��x���m��B\��_��쨽�;��t����e�3qyM��)ͨ`lI�QN�8��#L��<r�k�n�ȃz5APS�j �K5�[z��Fϛ���݉��@jv���+��Yeh��=3@�������a����jF�g��2�+q�*g���Iw��Z�/�M�)Յ���6դyC!��'��%k����(���8�Ƚ*Zt�Փ||�MS}t+������=��FW��p���$�^?�śŻ�)��s��x�y����e��|_x7�U���yܜv=:G)�~�p)�[��Na�u��l>
rH�{GTt�bq��׫���7R���n�	�ܟ"��?��f�̝A`|�F���L	����v�#xA4�XsgE ����;�6������0ȥ`�{�������Ƽ�&�H��y6H�a���`�~�F^��sf�jد749b5��pL�ӱ�J|y���Xԭ+1Ӣ�� ���a����m�mQ1ǖv}-;'�GO���#�P���i�Jp��gI�98D��$���h1���~�����\��)� �F���Ҿ&Q-�p��OH��H����n�x�%S	�ΎPpHs�T��?>��1&��2`��,�q���b���mK+
t�vS��}U�E�"��+1EX�-�3A1�LT�����G&{�@�%�GW�b�LzU���<zGM0��Fp3`��G	�&?OcH���C��6���E>�t)4SN{���r�dH�[Aړ���4:g�MjX�W��*=�0M@�M'�mHճ�`�Y���m�x�\�H�A9ū���a�0�Y���𞆲1;z��4�J��s��� ֘�=T�-�SE��#��%Z��7G���t[�/�4Q$=������Ɇ�M��L��>/���Ar������졏h�i-�K�;�lEe�c
�ْ̺��gi'_҇Z��{c@�� 'T�#`Ľ�,� ;p���a�8�-(Vv�b�i�}|�\s�r�V18����h�O�d��w����R��Sh����v���E՗���Ñ������-v����;)|�q�=G�ʔ��S�f8D���XN$��Ը������ِF�bC1׵(�!x!$�#.�C�|�zDN���I{g��yE�h���W��ȟ�!k8�u�q������o)kp�2��JX��k��*��>����M����w��Dl㞶�<@|�Q;��T�4�m�k`\��y����m����֔��yu`$��>��uiJ�4��<���@\˓��F�#�z�iĜc��˴�k�$$%2`�~�g����X.Vn���O}FX\����������^D��v�{b�Tߨ��r��:��֋��7��Kםo&,������m���fJ�R�H���ƾ��3\��9����l���	C� Ko��
*�+z����q���"�V搩�K
�a�U���@N�����3�	��P�h���al�E���odDx�y慪W�z'(�Ȧ��<�����x�YN�v#�'ȝ�,Hzި�'f+�jw	=�yy� �r�5L��J� D2:tӀV	z�f��X[q��5�>��q�0�C�ϚZY���3p��S���꾞��%y̦��C�}'�Z�v�!I�{��GQ����zw�<�r��UR츷q���f��ۧ���g���������;��@	��m����jʹ�,�9Ǩ1(�{�\�ᵠ��QOA����_u�PY94N�}��b�:-
*W��ϩ�.y�t�'	l����%�f��s�$i�@@��ζ�q$�?���d"R���E6X��-���Y���:�_Y��e�(�Ĥ�5��HQ��R���?.�0��CQ����Y��w���k

�����^�p� �n�S�9w��X���J�)J`�\oǩm�L�q�� b����Պ� ���e�yo�J-~I�]�D���M���y�IŌI�6o��U7P�τ�a�)y�F ,<M��1-8]YvJ*�.(&���ދ]L��`G=��p��N_�^�$o�a=.���O.8<!M�ܿ�wV�:lG~�?�s��$� �]L�9 #M���tЊ���)��ܒ�(q��M�����ǈ�Z�_2�6��Z����	m&���0H��zhi@�F�%���"��R��t�*��ɝ��G�{Ea(��\:r��r��6�˝Uh�02���"u7B1EZ��z��/�$�n/��pO�̈�dt�T�kb\1��3���,��J�(y������N�98�G5I":�(mM�e��Q5���@3�<��H����/:;o"?h�)����������q?��y��1CE<ޒL{o�+5w�s��i�~�W.���Q������B�K���o/@�E�Y���5n��@¹�v�ڽ�e�6O����=+�,KE���f�Z���)�yb��fC���|ae����m�&�t�͟�@��W����TWf�1��_�p
\>��1���o1zt�`��?e��Y�=���-��u�R�' {�$�)Y:և𸍉滌�+�ĝ1y��q>�pa(���bH�a����V�j���F-PP�1����w�3�s_{*��]UU�n'���%��xĥl�/J)D�Y�7h��ib��x�#I������_���<ĝt��ϙ��5.�X젡ǧ{�(�}DM�i�tAZ��F��X$�0�"�����D�{�qx���&�]%�J����3�\�͛��m@�����w��)�Ti-g}/�&��Ѳ��4	ƻ�S1"�v��s��df��1��6z-�����Ń�X;Dz�L4@]�L�X5��Ct���T\��]m�Q�I��J;b�þ9F�����V,1�e�<-�p�^k�?��td	�.Md!�p�rD$V'/+��ϖ�y!�?ֹe �(%�]7r��ӷ)>��MI��[rŵ��6k�$��1�x��'j�� mI�s���Ǭ������/]?���ĥ�Ԗ�Q�������?���������g��-��b_ ��\�������M�%��w7���8G�a"��z���W=�:a�~�0��8��q*;+E>���*�ĺ.��dÚ�xܸ|���G�Q�d..)�Ǵ>�z��t �9YZi�,?dx������x��O=����i����{���9����D��x_o�k
m���Q��Y�"h�'0�B�]��b�!�*�Xa�:geY�����y*�$�C�q�.U2ø%�׀0
[�4{`� o[=�\j1��������S���A�F�$���YW;@y��[�n<Fj��[V3D�_�5�'��G ���^,�ny-zXx��.�ʤ�+�=�@m�'��B)�W��j�6�2b�R�I�E}Y||��?�iX���J��œ{��M�1��[4��A�˛�L�#����W.$�iK0�3��>��������	ʖ&��fJ�|�I���=��{����9H��e��X�h$ԁ�O��}C]���:Vn�(\�0�n��#<FI�3'"|t�Y�1J�kK��y�SEU؛5�1���}�����7P�w���ޑ;�p�3����d���O+U���m����=0Ă@})�]%M�R�<܇����T^���@D�3r�� dӨ�W��lPA��Q�_d�t�TGx����4[s�ͮ�8�D*;�'���)��l��3���rl/�Q_�V����b)^��ڟ�o����ܿ�)���sv���CTEȨ��h�!`� KA#�XG��)�7��;\��^�lo%���޻��Y��B�˥��a��p�A����_[]�l楬X�2�(���&{P�����&+��˼��7�K�fk�?5�G�ߜ���>����j��\�^�AKT���J�����@�@�C�Q�zi����(\�	���kҍ�
��cfC�;D�k�Xø�$#����˕�~���Xr��1U�>�)C�P�}�|2I[���+,���c�6�7�{������Ԙ�rn�A���lRz�M�faad݇+l�6k��-�L��(ޢo�#t5��^��LAgma�t<i�{�"Ĳ8�J�P^'�=�����0s�c�4a����Cް1�PZo�} iB�I������턜5�� �8t�o�}���M���{ Hj��آYG: oR���
И�]��aU���d���E'�_�y�@o����I��6�i�2fȖ�޲ N�$�K��\�J.�����(��k1B�x���چP�L�G��?1quf�5'Q'(�v�Q�����w৹�^���Y~�3m� J����X� ��-�ez�߯���H��J}���<��y�*!�k����U������˷x�5˗C�Q�~j�՛�M�)�V�ǈ(ۜ�?�B~������Y9�	��V�9v�m���a��iН�����a��`FXc�|�<h䢨�����53�}�9FT��a�kzuS-˦LE��d��}�0�F�G����֭����Xm N�W�I�j���q�|��R�A-s������(����If�k�8���į�
	2��\� �)Ѭ�Ԛ��m*r��#V���)�?�d���I,Cw����.!M�jR�2���j<���Bfr��G��G�jz?�M�#x�-���J`��ƿfx�p�� h�O��0�#�w��۠J1N���)')~��%�T�{�|w�=�魽&�K}��k[���Y�V.׌�.������H�pti�%XZ�,]����&�[R߮��q2��䦦��Z�S�N �xNE�� nƣ�7n:�N��=�h�>87����W�КL�B,������Z�a�Fy*�w�_��Lz�Q����8�7K#
���� �.��yVQnY��r�wISDa�vF��P�Lt����|�N��. ��z]*�c�Ѵ���A��a���`Si��ad<�U�\'9�w9nm���H/�Cu
4u�"�>�Iw#L��)1��I��D0I���q3��/y�U��U^p�1i��J�
c�6q%1�ʺ�EW?�P�!p�p핅�shA2���y�u��Ѽ~,��Bnp�5:��wf�:�g<��;!��UMx����\«$���Vg����4kq⺷��^��t���v>��guQX����nW��٧m���o��ipN���|��a�F}.�W�(�P��<������?��/0�_3��>�a7T��{S�Ud�'1�D�E�ޫ֤׌g�@0��7��XcR� ��W���y��g֨ �G)���p�jӮq�es�l�o��(�*�+�'��E_q��Bm����Ex�F�F='��1��e��e�_Db��˹���;�<р�t�Em1�sSO��&��ކ`ca�ﾰ��sSL�6�J� �qH�x�7(����(_	��H� ^L�����xHۡ�G@��E�9�cc�V�[B��<#����x���(���ܨ�H����S��Y\��dSx���R	����H�D��/�KZ$)6^n�	tl�!bfF?��6�$�`!�Bn^K��������0Dkڵf�Q�ٴ���(o��[��g,���=��s��\淗h�I1ް{�:?�F��Mv�������4����C���,Y�}��t�Tn!�]F6��ԡ�	&I�X�E�������C�D�j+?+�m�NZR��L��*!׉v�y)kf�'�z��aX!+\�F���)bR��^XJ9;�=��7� ����"�,���Y��8����'�{���;�b軡�k��U�U�.�p#�q�m�gt{~��^^�=�`=�-�a

�~�-VM�6�9��[ �j5ˡ�CiD�~r]@Ҁ�iwYm��v�?h92zNr�#�Q�B�ee��v��I��_�Iu�Do�aKObaԷ�WA}>E���?�Lž�ۑ�޴�{̍��-����~��[3*�|_�w�Y�Jl�RƳ�4+��1�W��]s�W�G��
"&���p��1�=��+ݷ"�3�،�3X�`��Ѝଫ?��w}�s���:h�m2:�Cr�2i��8U�wz
bmx�%^�X�w
��I�M���B�d���n�V�4�	�4z/��H���o��p�*��{٫�/�
L��A�(�vԷ��*���{�rOUBkyiG�@�>���O�*3܂����g��Z��K������A��dS(����}�P�7���6���W.%��\F�>��j�v��� K9�n�0�aR� �K�'	c;�x�r��l6K��ЋA��%�Ȅ��Voh>lr s��69����t`�k3�:\����E�.k��G�2P�̀!��l��}?>�=[��2�� +�Y���MEڶm��ms�Ü���3�����Z��S-��_K�C�� {�H,̡p�_ˀ.���:s�$�{��������B&!�����:Ͼ2��ބF�"2�Zf�O�ky3�/m����R���ތ�!�I�i˾,c�J�#������A��ȃf�y�?	N_%����1�x�jk&�S�4of"DѝV"��c��ӣO��Z%}MNc�!y�� �N*�y���to�q����w~	�2��6�D���չ�yg�Hf>k�Q����*"g���zLFo�Q��:��7�P�?��޵e{��ø?��k�Ƕ3k��9!H�^t� ��[}-("4$�C4�R� ��>�QX��mɅ���u�|��#�y}o�F�l'^�o�g��1P�%4 7O��J�ؼ��,3L���j,�����B̗� n��4���H�&�E�-�L���K��K����A�S�����f"���ֵ�LFr�"�h�m����L�&�<�Z������1�8̈́Q7	�"{�2�O/���)�m�ab���%��)����5��ʨHi���ӷ��G��9Y?5@8���ذ�a������T�KE�k?�IR�����~�a�<����<Ut�a?ZW_�_��D.î.^�m\������2L�Я�rS��d��H���K:��P���SZ@b�g�#��gj������?���h]��%i� ��m�����p��8Ȓ���@�.SA��~&� ���Xp�e	��b�~��չJ52�A+�%T]�YSq���x4�cˍ�7k@����c�Z�)�2)����	3-��K�"�=�U���I�:�t�j<���oןu�D��,>�	�N�-)��P�[�C����0.�+]ۈ�J�y¡@�G�U�xiecǝ�a��j��� �K��?��TK)��Z6�&2��i��G8��й��=5���~�/���z�,H)'*��}���<k���~��ΐc�Fbߍ*}���� ��}��Q�T�($q*+��Qx�<l͛x�G
]:Fjݐ\<�n�c�4�8xt/f�hӇV8܁Q���s�W�O�Q/��xyc������W}_��3�k,v|a�����6s�c� ��j�E��ܘ�B�̇�HP��*qr�M�����������5M?�>;��}4�.TE�c%GB�3r;�,�.,��qt��n(�_-6��W��2�`9f��@�0�5]���K�M>�q�da���!�}� P���r���1��N��E�U�T(|���S�z�0Fm���zWË�_).���Nx�	�ߩG� �N_���#�	�$5�lN����O��~�cBQ��߾��WГB_��^6��b��$c�GtmS��	+���PŧF�_��)Ս�۷~��1�2��+jS�l�����7[>�BJ�u%d�4��*�h�K1�*�q�C�[��\'W�X�S�����R�X�Q�	Ny;p��2'@�T5f2�P�b��B�{��׿bѻ� BZ��Q�J�ɢH��D
S��}.D_N�T3�E1��=��)����*�&�����*8 ۼz�J���&��`��;����a�s���"�	���a��.��錦&!�T��z�aT��Y_��7�M^�zI3�� m����"���
�w1�z��|����>;B�4�\w�5�t&<r~��"M=�ǦHj(�'��3G�S�c���ڷYZ�ó��49������Y�rh{�ش�E�
�Z�*(�|��/ޖ2�Q�M�2���f.��lÉg��;w���o�¯��g���:�M㡣h�!�y���0�?έm��Q�M�����|��(��~���;ÿ��L�@� �����i�ݳ�D^ڧ231A{o&h#�9E��+tj�cJ�PN=�����q� ��'� `.L�ם���?c�#A�Et�Cô.���YzD�%w����� ߈���!���ࡠx�A���~��V	����G�	gT�Ѷs�6uŅ��E�g�d��W2���*O-;qeE��7T�Zb���-���_~4�U��5�:�O��]�6����3�!�(d/Y5��J%��/�о<��@г�6���ײ5�hȰ��^�j�)}�7OjQ_q<E��� �m	�`�D�O�k��iv׎(zu4�&>���E��,x�?&i:Ap)�sU;����[��:�e�����O���jcj_Z�l��T�#������/�;NR_��sy�&� '��z�y$u�p�c�	Od�� �3濴��E#Xl\C��8�r�3���Q�69y@����nS*�l���\+�����4�w,��5�1��x�\���v��GS�e�++[j����2���1������@��}i������	qv�!��g����A���FuW$���R&ZcW�Ll�\E��_q0�H�=�k�B��+7�X�&cB￴JqQcC痫������x�z���o�C64[!�g�N���t]�������3`t����6���}��\`*����62w�V̥�y}k��5*�����X{���������`l�M���}�PB��H���y�F���^{�B��ϥT�&�M�]b-�*�|�}\��7.abFq4ƇN\}֋�<'�Ar�����~Qw=����B7f%���	ͪX_m���'k������ �5p��'�k�%��fp��N�qkڋ��d��,V���4���DPy��i� �_:�t&��	��}~�X�<��O�㡠ƣl&3�'���Y����4wx�tm��X�$�_H
,�_�`��f2j,*�s t���]}|�*I�SYJ>�@��VF�ѿ�hc]��ɪԽnEgx�$�֔߿�vfc��̧uZ
�"����t.�����"���,��Ut˰ :�D:���8�jE�xT,�
^�fJ=T��|u��0�&�tr�tG=P�C��YWX�� ]�f���!��Qm�o��םv|�E0�ƍS:���O0"��E3����ΉG�5�̃h�:,4��*�����d �ߔ�쫺]ʲuDO/!Y���Y=�?�K�wl��`�N�f&��ܫF|�i Zޙ�/ϛ�4�*Q�v�8S�$��t���_����WX�+�Д��9X����p1�3����(1�~(�+�iO%H��a,E���~(���,"|VU	�!��=d!��G3Z���a��*�P� ܰ�~]��a�����:��a7U��{��6䐂�c�b�AѴ@�����m���y��i@%�l�݂��F7/��Pm��Ƣb�G���a5TyK�Y���=�J�A�;�X��nQ|�'s�Hp%]�d3Ą��pA�«0K��{)6��g�,���n������	�*��u��1 ˉ�l���k��(�p�� n-[���-��
�t��FmaR���)��xkg����!��&���Ў�=cx�By'�
���A�F v-���& ��h`=�C7���GS:�Ϲ�t�?�su(�n�G�������2 j���I���[�X3t~���ȵ;Yuf�-�k�((����k��s�vL�_;���t+Kĉd�X�gZR�=0����;@`�s[�ϰq:e/p��A��i���G�WO�`�k礮f`�L�x������E����U=@��^(��$Se�j�a�M�~D=�X�2�B�.��X�EZO��sp�@hʽ��u��b����6Bl��Y�����]��L����D��o��zV�d���� zs�}�zp����P�"�������F����Ҷ��(��z%T_�!,,�=�+���k�S���b~1��I��)~�7�J��ev#���۬j�X"�qB�pPW��6��k+,Q0���2Y��`������R��H����͸mIO��܆��	Ҋw�w�:�$/⳷���H���W_��J�0�<�,��wð{�F��������馝�%)b2o:↪�:k��T4���+��BD�֐�*���u>I	P�̗kVĪh�i�$�t��[�L-I��h)��oTF�4H�����W�����q�p��K� �c����	�󜬀�ls�w��n��}?� �M@��ߜ��~ti�S�WE��C�-��ɴE���em��u-}q�E�:q��'�+��d����F�[�{q���"3��;I���UÃ�x�mH�=����0��ʐ�n7���r�N[��Ҧq8�0�ޠP!G��ٮ���G�J� �d$�2�[n:� V�SǍb����r4��Zu'ñd^�u����8\Y��}݁R�p��^�7��郍�?]TL��������j3�����2X�@��rm�O�,&X����.6]�HQZ�@��v!lɊ�8��\]�]��Z�!�$&�vg�]]��E��]����|,�<v�����i�">�4S�֝W��ڳ�[����Bع�ᐺ�C��̇;Ba�V/���d�
���i뺳���\�5���&x�Q�v�`xj�2�%P:�z'�1e�r�� ���q�k>�A��$e�T*��˪� �5q/k����v�����nhg��wo��&S�,�����;��=M:���m1[��/jj�д�Ϸ�^r������ta;��Qܮ����7_q^�� �D�����i�v�]G�ƈ���e���!a�*68y�.�[텗����7V2�ܘ4�fn��|4����k5��(��+i ]D; Ǣ려ںZ� #�]�e�M7����9�̺`�]�&��\��^��D�u�Ԉ����g���;c	4�1�p���5��=\��
8�Е��#�W�������HAAR-(�[e��%�Ұ�=>���F��Qf�E��fw��SF]Ĝ#�������}�{�F�V����d[L�q�V�P�үz��E�|�����O{E���X�~��X�i�
i�
�}�0�)����n1=�w|���*������7ݬV�B(ā��G��J)��H���f�;{s��`s��P�%�Oq�����z������t�{VM�Ǟv��u9'J37z���!�����Ң��|s�pCI�1*���lh-bϩa��P3>����Q./0�2u�ʹ�͙��X}�K�F��
�CM=ү�;��x�R�P:����q��I2^	{^H��&�Ǖ��4]��.��J�H�Q��֪\��e�"���.׷$�x|.�]"������e����0#_��5:ꏶYgZZ����#�	�+�N{���8�z�C��Tb�A��[`�+��㎫�G��^
���a�c�[��I�����I��L�vxLI0��zJ��a�9�*��䳤
�f��|o� XW�!���)�~�؏�;&xb ���3Ͷ5'��_] �������w��D�v&��^9�P/(�\x�*�"����YN��(9 �	����$�â�V�y>�{�lp;F���J.��׾Q�%�Ɍ�Zj�\�Ol.�ՠ����eOR%��ĲdX#Ej���v�vh0�6#�Q��.>^'���S���i��Y#�������QS�٠��뎻3	�`����#{mhmU��A1$Ӷ˴��H%��-�Qn><#���ūI�%��I���z�a��?�k	���t������}�C`!�!���sJ>�^�B;�0���$.M�
��qR�F0�`�Y)x���u�	kih8b��zR��~P�H�kI���x��6�+SQBo>��e>r�]���3��j�gY;j=�|�%`��T�`b����Nw@�@y�6�jL��];�F~:��������L�=�%��1�3�ܿ"���W��d�Tj��Y�p�n^��:߻KĂ������ա��׾�je
U��Oꁓ4�9Mg9�eܑ�[��Vɯ�L"������~,C\���4�������Ð�q��l�Ɉ��OQ�R��fr���EXQ~o�H���(���y���oV� �_$�1��GKIv���By�d������N�&S.���H�����m�|��������;�OUA���AjS�p^�μ-R,�B�(/�̑j&�HJ�=��U��գ�55�2J�����`�P�ih�Yv+�g���_�V�s���#�/�걶)��,����S3ƫ��w��Y �"�L����!y�J}��� �l4����Јz�17�u��JB>d:����Z��c�'!L���aI��S�/�g�*�g���`]��-�<��/4�?��%P�W ��Qٰ�5݌����XNK#�l�:p���)_��%��A�����p��f�:��\�h�� 4�^؏�s	��_ūx���g�
d����dT�Bm�IALg��<Gy��⏯Ȭe9Tq�Q@Wc��c�V���Й�8�Yt�$Y�۹G]c>n�u�Z;ꐙ���m��o*5�} o/���H[�zR��t�gGk�!��g\\�K��X'�i�,�O�q��՘2�JXS)���gQ*�<�M��� �D-���CjP����صM 9y�7�W��g�.�E���_��*��Bn��[i%�v��M����h�쑅��j�\��4�p�n.��'�����3�w��SgO���ZX��d��
�d�!V�1tD+N!%F���pջ��*��b�4*Nh��(̽���4���-������Pǖ(����L�(�#7�2F�Yү���uoE�u}�{��'�@�q��FN��C=�$��і �Z��@�P��U���)��~�儻{��	˱��)�+AĻ��=�D�]������Ttl�w����-0��
����wտa�Uc4:zQ��}~7L�/��N:��t����@n��p�����V�'h��ya¹a5�3�|���~�cD��y�Z�А�?
U+��X�&�Ԩ���~�����0��2�ء�R�K��;�`̾ӝu��;f�#5�`�v ����4�Y_��$������Q4�FKC�b"LJ,Dj{��I�"�����S�
���2g�������(Od����~�����w�R�"f�����$#�:�dm�s	��f���cј>�P֝p��5ZL;F�}@�A�BH��@�N�Ø�w�<�S��"ؒ�;��e	���>::7��d���2�Yޑ���N�Hg��p	lDkalv���D `�^�y�<���m���ۀ\������p�g�������5'���1V�������A֞TzGy^!iU�af~�&3�p]�Q�EL�����{{��'��?�����l{���3>1��?^��!�-0�����l�Л�N"iT�x��A2~�F)�D�k�9،�)*4j���(��TCR�w��kAk��y�Զ*�!rZ��8���{dQ�����`N�@Q%�v�r���W�!��_ġ�17E�S��d7 �50�,v�f?g��t�W��~X���j��dr[�V�lJپ:˨��h5���=c[^r	�U$��{��o>kn���x�IO�H.�Sn�ڟ��!�I�����g1�:4hb��KV�y��[�4��6Ԇu/ړ6DǼ��<�R@Č)�=�(�0�W6]�9��xK �0A��U
�҃ /ކ�%�H����-X�MlRJO�k�-$Hy�6/��ѽ��u{%!ΉMS���[���__N���kNՉ�X8�HgB�` ����D�-�4 �3���{g(�+ ���;�_����U�|�5�+�Te��ף{<�!Yu��t�|8_ �w�E�eĩYS�~<.���Uw�1J�-��c#0T�!)���l��y�[F�-���N8�ԧ�u�Cp��X
�JZ�<d�����&�}�k����j\�:XP���wx�Ԙ�����׼Db�
���`�-���v�f^j�K��1���c.OI��gf��5�T�;ޜ(��v��5���W�2��� �`��M �'�h�|�1l�Y0L��l��j��B�B��Z����m���{2��%�J���w8:Z�����B)pKw  �!�4+�����Q�u���d��bW����9�TN����l}ώC���h�{�P�{� ��p�q��3y�U�)��U�Z��.�ܨ���)����X��
,��`Є�q8�O�t����<�TBs��6�Y������'+��T���&����&���`���-t�h[3��񼥟9n1\d�Ш�_}a4a���;��O�%��ղ���L����Y��I��g3�`c%���ŋxB)�y�˳�|�k�HuHmM�'��D�T.]�����q^�]u�߇Q]ď�E��aA]��PV�r��l����-�K�}������x�
q��D��-�ޞu�@|}�$�:H;�C���\�q�y���c�M�tŘ�=6h����\:���Y��ܲ�4m�n�ҡ�3�g�Ad�_�R�~���b*�o�)�JW�c�ֆ\� �g��2���F~�R�c����.�H��Vy<��΂UK@���@�>X�ty�LSA�COHŖC�`v �Wm߫|��nH�� �1�p�a�����\#��kp� ��`�2�K��1�إ��׳��Zx�u!O)[�׶`h�����"�j�Ȅ{K������0����&Y}�[�Ze�FY�h66rtr�K�O������*�H�A�Գ���	�aH�����k듢
lm]u�����<K)a����o '�F5��2�ϙ�>�<�Dn�V����� �dT�/�;n~u05����iEXT�:yb�7"i�/a�dO kfn��V����R��]M�h�M��C��߽�?��&��z�֊`tD73�Q���K*;���y��ƴ�oE'4Uǹ�Z�3L��h��d���jYa��i0g��w�mZ�X�|T�[pѣT����ma����*lp�T��,���J�*.%q���`E�n���'v2Ʃ/��J����cC����� �_��{�P�CC�/�`}{M1cD�1^[w=�!X��̫*�K6D����3_��?�*�'�ɬw�CT���C-b�1-=�a��D���G���s�u.{������#O�g���#P{a��M��#jye�h5�tV�A�m��U`J^��Jx�Z�T[�Q����� �dpHn�_F�|8Ы���1��] ���r,`Gz�K|��� Moj%�����o����0 3LvN�|E�;8�ܛ��FdC}�Z�EZz��������V�a��jN��?��̏A �^2dvX|��q��NtE����d����	qgXן:��,mAWiΤ�F#L�E(��ߢ[��=z/��r}��'l���c�"�����w����0I����PN�9X���pw5�:�h��cU9����-�5�#ـ5�k_�5����8��{E/�������KM/2��.D,+�˜�I���v\��3��T����\AE�վT��5�8���2v>�xR�lہ ��x�Gd[9�M(�?��6��~�(��.��!S�R�I�(�*�@D�l�dn�_��� �@�-�Y�un<M��\�(~ד��t������04"���S
����Y��������3�z��>ՔaٛCaߤ�1���K��ˀ�9о�.��Ђ��i<�3��hk<5�l�q^�� z�.6�>z���k�B����zL�:���+5��q�H����:#��o&o�z�;~O�F�?��A�#�戕�3(V�U� 
o�n��I?�!�@�F�f]*Cl��1�G���Ea]��n��o��G���,f#E��e�E���&���P������J�Q��&��_���*�YH�H8��B � 7匿�W3�Q��1�QS����r���ի=�KG\Yg�o�u�f5�eJ���]��	�p���Ĉ�i%3�L�YHZGn�q��`����>vp]8i�R�G�Tg,��l�� ����N!�8����}(����K�߰��{u� ��d�jT)^���x|�l{c�ޮ���(����l][,$d���'Y��V��b��f��Z�棠V4�)�����yۘ�y��e=�܍��F }<% m�b�y�R_7@�Ԩa/d�_Jp\]�"�#[���?��AY�-+�.m	������!�)��9TrP`gW�w�v�/1����J�D~�z�PP�D������Vn��Pbf�XM�_0EZd7��s��U6�8̍��n�z,4��j<6s�����[��:��r��6��6�!�6�2�n�A>��*̻e�U��\]�%�Q���p��a\:$dY�6Y�(x�b!C�4z"�j���G�M-���I`R���bH_�w��4	XyL�@v���/{��h��@����D�\���_N��pY�6���rx�Ϗ�H�	��.W���V"�H�K9@&
����ώ�)�KMέ�H[)�<I� ��;a)��O6�Z�1�J�\������>`4��}��h�wPۮ�j�B��n�v��4�!&�5�}ZU������
�'.����I�ss�ȵX����'��Ԟ)��}�����O?���{o�9���"�eg�I������5�O i� ��u獯�Ǌ��"z�p�n烧��g���j������?��l_T5���D%ָ����5aQ���"���:N���ۉ��r-5ܱ��_��}d��������To�E�\�aB�ZW��װb$��@D�l�/��xh�_��0b�5�2�x����[�J������4ӗ�k�Ԙ���C�ւ�j)�����|e"���eB*�+8'�5?��T���o���X��u�X��Z&"��Z1�طUo�S�
<��|��
�J-�b)��)�5� Ey�J[>�Ҭ�'5�s�R������$;����Gm�qM��}u��2U�f�t�m�+�tyu��ƌ,���,V�5k�R(4���WBu�y U'���D�Q�00��d������9+k�+u���U������:6�����}�b�Ky�~�;�ݩ՞O������/��;����'�]���<~v.�Y�##�� 5x�0��aY�݊�w+JT�֘�e�kt�j��j�ofP�uL`��0�>6�@>�aO�G:e����@���<I�ыI�Кţs���-6��N,�N�����Ec�֮���ON�#-�dG��O��}
.��rU��}�s�`4�0Ȝc^�Ńq��=���ïA�v�	�7�zW��/�gc`���8:����w��2��܊��&����Mt���º.��FC�=i�o�����pKCʱ�ѝ�1;�UA��M>�����F�pX�qG7����R�0wU��m�ݚ7d�瓝Y%�#S��ߤ����*$�g�K�z��K�[��	�p՗։=BF�PML6z��ȹ�<�P ̯���E"�=��aX��\�1�a�+,��,B� ����)T��kN1���+`��n�k|���2?7.�������a���F��3��Nan��[_1Ch��j��}7=Q��pi��������DL�8n6̐���x:_�rZ���#l�
Cm&]�=�7ŭr��6�p��d���~�lU��7�,�(5?fc�|C�2�[ځ�-x��.��R��"���+?c�X���N8P��1DW������T�B`�̝6�W�NBQm=o�����M�[��s�'p�<<,����������Tk8F,C��ȡ"��*b���/*���{MRH\�!�PT�GI��K"�a$�4�]vnJ��i���B�4bRe��/*Z*ݐ��6/�@��b���#�'�%<!13CTTt��$�-��_`��Q*zMH� �t ����sW���#Y�
_��n�/}��o�*�dø��5�)
-�����z�
����*�SQdNI���P��*��9��n���]j��/���A���	��D=ri~�`�co!'S"s÷6�w�H���㛌�5�pȃ�u��P�[k���us9�������ЪC�4�M��p�k�}�_�@���T��K��G<-p&hg����\�8�r��<��l�������?7M<ctDR��2�®y��.jL������dw��K�~w��	2�Y��[���<��g��l�8����G *�j�F���y)Ci]�U�"����j�M���j��2�	��f6~��Ie����Z��U8Ǖ"_�M��yF�'K�#�u|��~z*���F<��F�HI8|*A6K�ӳ2 �Te.?����&R�P.Q������a��C�xC��J�^/vZ�:ݳ[�~e��"б�{m��"���0��p2���LT���^ �M�tD���_y�� ���qޒ=��Ր�k(eN>M߈'n%�N,��6eڑ����V�)�VbW�X����0�5�di`�غ��A�ڕ%٣XE�Se3�-�����컡�k��Mmz�	��v����*>��M0Ceh,�Q?�\zn��#��Q��5)���[�Vf�1/x�)���KOz��[jПT?���k)J[/��K1c�\TC/�=*G؁�;��v�vX �. SZ��Zc��8�9U�0Z��y����1(����C�d �k�4�WZɝL�w��δ��CY��G�Q+�Բ-m��\���+�.豵�p�(/�]��0��y)3��%�օ�*4��IP]w�
����3��%�)�z�Vp.��ym̌��R޽D*�{���[(:�&(��+�TC5�a�}WI�)Ɍ=���MB8��ˮ���he[�ʹW��W9�F]�g��]�����wV̜Ia a(�y39����[R�5+���f�l݂,�$L�յ7.�H[}�nq�ӄk�W}���oQ_z��k�w]#�
ZJo�<%R�iQsU��qh�8���=�K�Mm�v�iΟ��u����{�2���}w�B�.��V'�m���
��� �ؚA�����~D��k�ɾ����;������Q���w-��h\AQ`�#�[tI*�Eay�/Z����2
���0�DwĻEԴ���q��f�ф��o�,hߞ����L{�CyZ�O�yWG�Ч�٫�Y��D����;�C"�II'n��k��C|d�B�_��L�%���"��q�h0�G��scy��Ϗ�I�H$�w����M�i���U��"����;��k9_�"�]��w�
���D������g�ui���V=������ᎌC5 +ny�Pa͸���]�H�a����)�� G������8���4}�à�ߒ�t�N���_c�tqI 0E����O��$^�^�=�O���(�eh��9#N���$�]Xj�ӉqG���@�Os'+8m�\/9ń9�t?Xo�9�q�~f�V���ve0�:��	�]�h�b�g�a̐^�����i��O�ɡw1�����(�u�yBu��$�^�	����X�����gI��S,�b;%M�	)7���&N#h� ��go�8�����V�y�S�QM_��h^:�'Er�H���8�p��V�̥�WN�5�9�I�N������U�[��࠲��ðs����͙��`ܨ��į�V�/S�?��g�����c�����yYS����y��,�-%�����7�\�r�!��3E���?Yu++1��F�� �r�苫R
�g���9�#}�Ȏ���$.oՐ��6�s�P�,H^�����!�[�VȾ�}l)�+�n;��nPk��,]��b�n��	lLS�_��p�bf�=�����dl,XKDbh"�U#9�F�jv��{ֿ$�뗓��!t�,�4����ї>�����
/�s�p#��*0A���:	}��<�ϛ&j���G(�����Zs�i(�2).��$ݡ9@ű�p"�_ڤ��5ߓ[�ፄp��՟��~\-MP3��߫���(l����9k���ap����'�FT��+�9�I���'�ZȪ���	��Ӭ���8���<g�o�8����!Ea���y|���r_
��zw�9]����Yr$�@�g�E�.��'g�]��ow=%��Q��FԴ��ii�o�Ũ2�Fy��YR�?6_����\s|�>�]^��)U�e�;/j��¯DG�~T��%�o��W5e-0G�K���`�[z���#͵���Y/N+"��	��,`�����C�Fo�Vv>���Z9�/�"�a=a+^�D��F���6��8�qg��e�0�a�mZJ@�+�����R���m�,�<<��/$�̣ȉ%m�6" ����S@+N��q�M^x��^��c;:rcB�o_�ā��%F�V��V���3w9:H����}@T"�Gnb:J�m���a��W0��@u��L6�P����r��r�qCk�%�X���:S�UZ�kB�5ٶ�=Gw���)*݅�� eDiw`��3�[��u��( �j��Y�h#w��2(�Y@a���Q��� ,�* ��^u�V�d�H�,ⶔ?���Q���{=N��Y\���4��ƿ��	���d�څuhRQ�c��w�4��:O|��N��3Q�����hL�����"�ȞESF
FX��y�\-Ƣ�(�`p�~�d���d��O
�j`��E�~!O���^��@L�bh2\�F, ��*��7�P8�gjV�T��Sǿa#=$+�_M����㽞�ǡ��o��D�es�q=-���e1 ]��/qޡ%~�Ɛr'>D�ҡ�1ۻ��EO�9���V����9� �y�H'���	#*լ�8�N&I��;S�jCC��fW�!I��zi��$�����+3J�'�ȑ6�{��L6��:�~>�ްS�/#� ͉hޫGd��(@#h�;��amGz�H���p�T�0/f��ֈ!��!O�CV'�L����$�a�Q>��#޹2�e���$$��C2;���r=Q��J�y)�*Ew�֛S���̈́Tmo@��Ɋ����Y� 7��OZ��U�Scڮ���;��M;�q��mg� ��E�E��d|�X�����­>�\W�6�4��EJAwE���d�p�{��@k�/��A8���|Ǘ�ςMZ�io,�r��m�����x'6��sl+ �a�mm_Yl��
˓fɇWq��+]�r�ˉ�̚I������l?y�_k*��0X�&��u�y��x� ���v9�W��u�#�fC�7L{�0p�0�/	\����P��f�;Ɏ��{֧��,�R�I�O�Y)�Y:P!�g�Jר�]2����)�d瞟Q��⟾��(��`d���r~%ߒ�Y��Y�g�"�st#P�O�LͶGV�>�>���f��VI�ڼ���,
}(�����P�֟Ryp�f�,��o��rw��SSޠO�ޓ�x�W����ٷq�	�1Y�<w�Y��H�2F�5�Ɛ������0����px%����Mq��h!>�g�\9�ߦ�,��.g-�(y��u
��LV��

t��֢3���ð��dD��eç�m�	�[�|l��a�1��k��	��� �h�����,��>w�����M��W�N $#�ױ|��F?M�yA���4 ��b^\���<ъ�Sږ�N��6����u�c����}/���<�t��m��ɢ������i0g:�J��E�}��qT�I��kԘ"��E�/����#�'��y5&��O�#����m�v�6Je�ܝ��b�B�_�
'�M��\�"(ü*��`?&���L�h���n���O|"�>�B�HMsqi �Ņ6M�a!>�c ��ؽ���E��ug����fK%7�}�E�� h�
��謌�{���ǚ�&��EC�q*�Z��|1Y�_�h[zg�o��vF�>},���I�?�<4+�%.�7w�zS�U!�i����9n��ӭ6Vh߯����$͛e6�7�_P)dv�QL4�O�(��	�IL|鼁t�Q;�����׮�mS�8��8F6F�O�E��S��� ֪9/�X���x��q̸��̻�|+�B��Ω�4c8t|�y��+�[���b,˼C�F����
��� ������I�N;�LHf��A|f��Vk�fX�t�������\�S*�B����b,.���=�a �D%]�M�/�9n�c�V捾� ڄs<�m~�pu����A�_˘kJ��²*ޚs��>*szȰ�[K��#UJތ��:���G_��嗓ې�����;r"LH���K����i�ig+��{�\�Oe�"��E�A�$������"�8�6S�DB�W��`�EԎ��`���F#��I�m�(���{��(����v��G�!�g������8��/.2�^�R�/nX~�'��M"�\��ⵜ���s�&Y��_���������9�'��Ȇ2�_C~�5��-&P�4��R-U��n�Wb��;����-s�A'���2BO�զ���l�k,�{m�p=���,��N}>��y�wu�EUy��?� (�A=��>���)�wL|��1����d��1��Y��S��������h������������I����[[i��c���s��%"��HM�q��F��r�ެ��f�#���5�����q#�v�9ۯU��� "�f�Y���ˆQ�֐�,v,�����̮�(ĸ ��?{YD�-����b��Cn�u|htPmPjo��������4|����á�<#��U��1;/B����b7�i�]D��0���\OÑ:��[�DG)��N暌�ߧ'�Q��j��ѝ�,5�P�n�CnT#�>r�s<ċuJ��|R�F.�2W�|z��$�3w���_�o	����X�-qb�c�0�n��a%A0|���nV!f�s���|��5�ԡ:���=:�p ք�f͕����4h�QA+wq��U����E�k��3,b�Ņ�~�t���|@V�	V��'�K_�D׆-�����0�����/*�$���A?��j����9� �*-�5#@�6���������O3�1���*�W�pSD�F�q\� ҫ漷W��i���~�0����:�CI]~�|smB��>��"���L��"�$��KzI�yl,z�V5b�<�Q|[L��ɛ�Ό���a�9����_��[_�M�v!/��@�iGL�J@��i�A^�>�ē��V{�>@7��\|+��"����hkꠝG�@ GRY�Ρ����f�����ZW���fGL�ъ?�i�&J<i�L��8)���޼�ª��՜�!�2�����;1f��両,-kq#��{�|��T����Z��v2歁�����{��Lpk������u@��p8$-gJXaECh�NFCL���:���:-d��ﾏ�@�蔅b��k����>"��\��@�fK>��W��*�m�U@��o�ʏfhbx�󝼱�%e$��';��K���a�^�mI=[�)��ݪ��O�"~�K��܁J=3gZq #���G���B�7��[�|Y��X�ih�ɗ��7<$d`����+��q͢u2fEr�����j*�1��t�/�%#Ig��b��,t�����"�gtx
ƀ���J2ā)�m�2��tlX�JtI�A�C�� ��w;��R���y�!.o燛+��w�Bt{��;2b_�L��C����Xnե����3�sƍK�1�D�4��֓�N�c3ϓ8��y����%6���up8�7}������~�.`1ԛT7S�[�'��^�i�v���>�Ѯ	k��q��Ol<�a����!��%/�W\5�w¾45Z�D�ȼ�2z��������f�%��n0�	���O���=pOu�PM#�ێR��
�@jmU�]����[��&��z�=u/t�Y 򳩬݋�,�(����v��\�;qA�6�T�͢���\Bj)��lT�a�Rsd	����F����P
�ƪM�Tv��q0�%���ʰxAˠ5�`�p���!��^K���Y�ځc9>�8��%�?A��/�SK0�xJ	Bw��._9���K5��t�!��]��q�WL�����g��2��J��{���L0����&3k'�l��|���D1,ߑr����O�8h�=��+8��R�� FҼ�]��v�ca��c�0ڴ��n�V��.~�3�7=�D�!�+sg�i���JB�|��Dw��i�7=��)oJ$�o��1��<�6�Z=�U��)�}��� T�l�b!���$������[�h� �֔�������M��a�M���W��Q�KK��@e�F9��r�JO��ܬ�J�vIç*%R\�>�+�E�ΣӲ|/�!��ix��3b���{���I����nZ��.Vn0�|ǉ'�����4�����D�/_�gw�6F���dMw��ࢴ�S��?���w3|�5w���"L�B�z!!���XK�dg?t�_�X�*�һ���NQ})�i#WT˓.�OC��o�R���'���o�yl�����yA_�V�*�j����Xx�"WWK���=I�J�]O�E甽^u�_�>��G䓐r��/4�Ň[;�����x�.�qP�Z�NɅl�K0#��U��Ժ�0�l�͂���4G���p�.T?�[	U��ea<��>w��^
��h�D��#����Ҥ9N�f�3�JG*{�Gӹ�qr�"��,�EE��U�~ci�uN3o�	�{(�f�K�="=���/Q�M
��=9jY��s��D��x ݜ�����,�Ҵ���v�G���]c{��)-�\q�Ā��a�>��{��Fp[�6T�VC3kHx!��MG0x�ؼDY��H�UN�HO��R���(�����:G�}dX�ͼp���4'
��%����L2����H��%�ϡe�Nn3��s��}tn�>������e@}��M�����(߂��Sh���f�+�������,ڰ���&��~\w��,S�DjN��V��V'Ox�/"2Y����
���*p���yJ�M.>E��A��!|{蟖n�h����܇�Z��@��،������
YnB��� ��-KU�5k�31��@�F��>|w��vT�}�XA(��i$$+�wt:o���?n��`�84f�#�؉c#B1�Վ��B�����&�7���^:���&�1�l4h�'"��f��m1�r���{&#YK�H�*�"!�l�������b��n�֊-�������7���y����Pf��66�6�×�~X�=��F�E��4&��\�N�?by酽r��8��t��[%�/��Hӷ�L��X��V4V'��&�@[�w��	J6�ѿS˿��Oܤ#<�Jhv�J�Ỡ¶��V\^T����M7�ΒIl�1.�1&6Ò�i��p���re$�����p���afWv�Q�+:_HA��YT��E�m󼥡d!���+�l!`�;�q���8I�?��C��ڬ.Ub@r�O%hj�!AŋT���DU^7{��}�k�z�챙$�7c(n�"���ǔ�ߤ,�"���<�n�yn�#0Ƿ��y�����w!�D��9� 5S�tn�PUADq�\!�y !�D`����Eh0:�����'ԷR�J����שVY!{�G�����K����ڙ~�Zm6��/�e�~��a�`��h�z1�Q��"��1�}¾/�T�ͯ3�O�_fxJ^�l�p6��Kѯ�[�1�
����6O�zݜ@�g�J�l�C`h~\����eu�1۔���d��g4��F��f���c^�g�I�G��ȱOS�9�.,�9t�c�k&���=��i�W�!�x32�m��`���:��W��y�y`-�+̖����Z�3�
�7��������{X����-v����Υ�]�M�S#9�7Y4�.�#�y��F�[F�lN��vZ�e3gJO�C{i�V��<9ie�Y�@Ū�JTKņ���\O��C�(h�jz̈�� 5�@ړV�S	�$(�B�U���]�e�I�.���U����߂reL� y�KZ@�u
1�v%��֞fl��=T�v����8<H�vA�Q�3�����5���r�c�|P�S�M�@��ڽ����=Ys.$�.�ºQ�����ݤ�g�V�����b��?z��YZ;J�}�B5Cm"<o��/���dPmt��骐 ��G���/�	e64/@wD4��_~؛:�g�7���m��\6��K�<�c������}� ��d�{+�qE��8=�z��<@�ͲK!�(�?O$AoU-2��,�O��7[��%���_�uQP9���~��O��(Ԑ�4�:Ԁ mE�M<�E��p�9T�`A�w���8�|	<�u�'M=�0��5�� v�(n�e�̭�LҀ:��Ie��7��:o�/!���C �:U����2�+$}[�����܌��4|��=�q	�"#`��?�=a�G!w���,�֖������t
Z�@2vk,�I� p� �n�����S1c�=���C+v���A�)���k�'QI�8�e,+s;~�6��ُ)�[w5�U2ϒ�a��>1�������;�=u�~{�AEVEj�.5�=��|K�r��[t������Iu��fJ���@Gl~6W�1mG�kƢ�^��$�!�}h��	p���u�l�����]ݿ���{N�0�6 >�j�ٸ,�U������g��� d���E�,�G�H�2)_^0�!�{G�ؗҠpy���A�v�'���D�Km��8��UOQ>�I����J)?^�1�!��{}oPLvn���ŧ`߱�+ 1���Z1�����~��T���bh
v����GW*�����c�F~�B�q����� a��R��"
ƽ�G�R�����Hݴ�5#��G&��p��N��a2Z_�l��68ه��pw�0����� �|��Y����z��Sn�>�ѦZ���Db�wrﳊ�R?|�R�&I͡.{E턌�F�fy��6��׸�ĩl>_kVYe-����U���cBj��фhԿ�S�i� ����d�]���֩��9k���KD�<�c������l�1\a<ث���T��}X֢���[V���T��Ի�����cPX�����۹w��w�ܑ�p�a��*�;��GB�R��x��0���S�o﵇u�V�����"�|�a����e��G!�+.�\��U&�>WY�"�y�0��6�z
�k���ƌ�P�ִ:���E�5,�j��*��T����wv�>�[�;��z�d��,�YB��V"��|����s<�3"`*[W�|�W�a$eE 0�7:�]�O�[�t$R�p� Rr��Y�S�4̣�%�m�!h���'�@Py0��Hz˕���e�*l���q�FE7�	�I:�$7+���)��X�RVI�)	��tnt5��p�[D �!�+Lȃ9�����FT��'���P.	|������h������n���W>9��ߕ�g[���fK<I�نv����%�y��^����`��N��N�ck��),Q�˦�>�"+̟)�-�n�I�Y<V��݆_�ԛ�ne�o�g~^M�&AJtVE_�={-D�W�]�� �0��3���I)�啶|����F��&��c����f�芗� �.�/!��.���9O�w���N�* �9����~
m܄��C!�
��2;��(BU���` �z�@F�ߚn�A��M�A=�������ۃ^��&qrnj���s������i��|b�S��+E�'���{��_Eb�ãP ]=��ng|n�gMt7:G�Ô�8y�^m��P�}F��@���n�G�<](��<\YJ{���c@!�q�������Llȴ'�-	/)�1��
ƀ�N)y�2��������[ �� n�
O���!��YKX.���lO�@z��-��ϼ���aB@>:�sr�}2�Ꚅ���5 	�_qE;��6�"��>��D٥+�Xr)h�8��6�ƕ`�1df���H�%���1��J��_�m���  �������n��A�rb��xU�j2_���W��(���m�A�O�BO��m~ȵ��	/���2���l 02�i���C���C�b���Ͳ����I��-����?U��9V���\51�Gƥ�����R��tc�h�bKK*&r��O���ЍN�g�>v~��f]c�ڵ=3π�r�P[�Ni�7��,�Um"�mݳ�m�$A3p��*'��xUA�Ԡ^�>����oQ��Mι�f.o�f�STW8~�n����7����>���)}p���0���5Xѿ#�n-"�R|rP���BMi��a[��W�q�d|���n� �]��x�t�)�l��������ag�|���'��%S�Ze���"�{�0��Iw}�[�[�-n4�� i&��⪖"�
��� T�kW)��T��0��I=ݘ�ܩ��u����v�Q���
��};ڱuusj������uo�$S� ���AZ�f�� �+X�JݶS�#�ʔ�p� �}@~�����&��z����Pj�1��S�U3�]D�C1�ᦖ_�f�p�[�)�|jE�>!��4��W�>��c8�t�s,��!r��1X+�����[/Y��h��q���1H'I9�gIN�|)�	�Y�΂	�$P�Sc��g���e�4���zO����xae���F���;��?�~�0M�6YW����o����\��H��G[�U��40c���c��_���C���e��E'��䱖���ޫ)��F&�z��z�(��;�,�R=�@��C����u�zq������}��8-��K7��S�d�R�u{����4 ��IAy�T}� x���Q�z�EzMoc7as��|%+�O�.& ]�V��8���G4J���Ͻ�KS�����)��4��[*�8�R��(Ypi�(}kj��'�I�O��N�d�)��rx=�O�TQ{?ن�x�!����_;�ƫ>Q���M{ ]�97B����H�d��i瘾�P'mq�@ZTS�dAr���sD�� �p'��N;�Z�/�Le0wJ�`(�|6���.֭�ɨe�SJ�
F�ϐ%S�Q*=�[���2��*M�8��k�]��c�-8Br�T�Q����K��lF��R��46���Q :Q��@�N���I+#�:S)6�x��t�<K�om��P?>�=����w=~�.�/�'�-6hw�I]�GJ�x2��� )Bېm�n'��ڐ�9�Z%���I�e�Xt�r��{x�២�ͬ߶���z"���`��k�k-�ߔ�N�~���xo����H �[�3����=��,��9�	4�1#���SƟ�n�K��рF;�� \���u��q+�s8���U�;�&q!�-�o�n"�=��+��
��?M=�GЁwl#���g%Þ�C>�����J�����[����;����������{#���^?t!��W/>S��Dh�p@L>�����Uoh+�4×zI.Jd�I�X1�G�a1-N���ES��/�L��Z0v=s��b�Iܥ�"�O�?��1#g=֐ ޣ��uV��G*u�a#X�
?Cre��6�j�:�/~::(	�9h�ww�y�L�������؄/2y�n>�H5�ܭ3.ߌ� \����^�J�ێ!�-�!��uBD1��}�c����!|�.�/4do59�q��駚�%=��tb���3~�!�1;��,��/miG;����D�X��!���W$�'��N��N���8��;6�1TO�O��%5�����Y}���'d�p�����oq�YN0��`�--!�g
C�ꅂ��
(�w@���h!ۂ�	s�S�l�ۑQ0!A�"�ؿ0����X ��s3��c�^9��[�u�lM�͑�p->2dE֌2��"�~�׫�%"��_��`�y�u��T�5:B�-�О}	 y-j�Ɯr%��\�y�C�D���A�4n�Z��@�HiV�f�<P���)�|/~^��躍@XrA;AI&t���6�2OOW�\���Er�� M�"b�w~��	��S�����E��嘔�̰VR��^�>B���c��fyDl�	4����\"w\�=�u�5��(���hԃ� ,mG�c&Z��%q�)�ʦM{ğ{-Ik��~V��=K��ɚ�UT7��[����Y��nP8��O���p�X?�#sR~�b�v��I�<�7��W(XԄ�����RU�Mm�,@�[�#4�� �G�h��/������ػ�ppu?�`#u&���C��� ���hgY�`�_!��>�:�1>�4��;���|�)��IUP~'�wR�N�S���}��k6g|z�Q�t��wPZ1V(�ڏ7yH�� (J��mO�3��t8�I����֛#��P5s�SO����}�� b�0��3i.�Ep�ԾdN�͉�A���}�c�\��$��\ݫ!��C(bYz�h®-����j�q�	R�y���@�7kp�-��J�����hmM�G�x�d�V��΀�Njq*.2�7�'3�5�t�'*��㮳;��8J(
�g~�#א� ����4�PŇ�*Y��ȝ�l�&y��Z"��M�W���^�]]5��9ߤ@��.�5G��l~�q�W����#N��ӛG����I�	�w<6�#S��0���3���Yk1pߕ���B�_���~�d(����7ܴ.\���m60�@]��4���R�B����@2Q���V�G-� iZ����G�2e`�Iݷ�M�z� ����Z9Ȁ�Uؾ�q2{�
h��e�-˴1�9Z����Y�(1��22y'�M�/y�Fe��{}����
�5Ơ6e���^"��4,;g��+��	cd8S�v��j��|��l���ӈ�����7��,W֘;t��Q�T���^*�H�sW�Tc`�>u@p�ߘGV�M���f��C&����٢wT8¯tռҮd��YZ��a�م��5�W���Lz�B7�_*{fN���Z��c��*R�J�Af�ڠYw�~=pvg�a$8e��� ����K'������^�u%*��G��G�X�]�%��XI�H�7b���d/(���=� E��x��$��
�[��%��`<����f�a��Qq���2��m��3�Jti(����O$�`��c��}����b�2��/~&��C?��H��H������z���چ�����P��M�Ӆ3d�'��Mi��~��_-]��EU���M���T$k���d��?���y��>���  �m0��s�\���'_��V3���'il"8���{��(��7��VD�ar,��-����� �m��KkPsD�?��jN׶�/@[3�7.���c��KT%���_Pvn'�r��9+�䃾okƒ�/����wkޱ�N�C?;@�r�^��({�t
�����q����3��Y�z�m�\�l�����g����*�}RV�t8���\H�iR��h�MB��l����U�pC�Qu&�c¥��������'y����^@ކ&�Z�Jx,$l~�K{��A�_7�ws=_[lsK�<-�f��7d;��1��tF�<�k�ޥ1�i,�Idl�ѱ����$�7�Ă�=f��|:�.�g8Q{Ӵ�}�͓L��N!�9��&�׃;�Vqc�.у���t_ Tg��M���I0ډ:�zB���a���<b:c�z^�5{p��=I,N�_�u�?�X޻���5D
�o�N��ͨ�fj���n 6�����Y��)r g�/���@?��5N�yH��x/��h��j�a+�[5U�n��`��
��K�cΪr��$��u�,��D0[����o���I��T�JS7d�t��#;�v4N�J����3GŽZs7�;�݃�[&����& t�RȁBY��=�t�*6�vLa=�/���y�w��9�I���%�+WN*���kשU�Β��-eI�O�?�걮(:�;ʼ0M����|/Ki'�E��'�*�k��{��]�����᎞D���Ϊ�}哎r�}��aa.\�>� �Yॾ����OR����Cj̘�^�j���;v���<�s��o��dRX���\B�r�)K''�ߖ�Lx���?Ɣ��	o<S�S�G�˙�& x�Tnxq=�*�?����׻D} ��Ȫ~���_���!�*��POu� �3S�#q��U��HWԁ�
��ԔoΓ|<t>�mȽg��QȢ�H�
��i�D�abZ�J��4��J��d���f�7ۦ�
�UO�s��j[n2��=J�u�s�Ê9a����>H���) ��9J�ϧ�¤�r�� P^��'B�-�E��鷃�r8�Il�+��z�Y����)_j�j��GF"?(��ֻ
{�8�����e����o(�s���;�j�i/�\,\�* 7Q��8(+
PH�شtY�����S�Iʥ*��Β�+ɛ�H��o2���p�m�@u3����Yiо�>Ȕ=�T;�{w������Xh�r���}z 9������7eБa@;���U�
�g����'�6��Za	7���b�B�~pT1�O��	Q�s��D5�	ݢl`{,����3\:����G�pR�����Aa;[yn�JЯT.��Q�n��Y���0W}�E~�*�;��@F���	��׀���NB�AӰ�c2�ݑ���UJ�����3xk'� ��;y����Sat�C䃌!����V�|� �����Z ����i=�qD�^!E�:�
"hx_ď�
�������y�9W�V�sZ�trkV�=4/��S��|�@�Zl�W�;�/�rt��8pcr�q(����$f5�A�[�����9D<}��������ܨq��j�6�z%��_���.�G\���|�����4#S�7k�t����!U?s�7�pQ������]�r�B]��wk�[Ӑڲ�́�P����a-���W��Q#�n�V��{��A��������}�\�\�k�dA�|=�\?����������f�o����iY	5�ۗ7w8��~ӏQg�=�%s���m]C<�����ۇ�a�3XQ)�	}qMP�K�� �tp��������.����:�����Rߡg�%U��&�^U�ߺ�0�/��|;Mt�M���\���}bh#� ;����p�:����%1��~�j?��<#/�'��y�(�i�� O�����"-��}G]n�`Y�v�h�DhD��ຢ���ҽ�r���w�⇯���T�i�shҲAw%�Q�e���w��Z��P�A���������v9>��8k=Crۤ\���$=�PH?mJb"��^W�+ �����������-����x�Ow����C�e�R���W����g#,�s�V
<�.�Հ�c��mŚ�������
�)	<��{�I73T �Y��Q��sn�s�w鞐{
=�~$p��̥@�	�i������Ao��VQ1�q�\?�\r|��f�1���F�A���<ڭ�Q^func[��{#,C� Pf�i0F��c����r7Bx3�8&y�N�d�ç�	��.Y���s]8�umY7ia��j�U��T�r}0��Vѯ^�C���p���m�'U����%�6J��mK6��3��&&*���Ù���>��<����a��bw|ϿA��-�1�<o��u_t2�I��|�F�#�}g��I���u�?�V�<K�8�����c�"Q��4����U.1)\��η�R���pM�g��OQ|j*�}��k��q��N��/Nf���G�0/K�;��{��\�3�kb�(���7���x�B�]�o�=��j(m"�/W��t���z��l>�rH���{�2�.�M�A�O�ʲh���!gW�;=^�u)=g�LL���Ө�G'�S���A�e>�_��M"��T�� ҝ�$#O�a�_�*n���1�	��o��|3���P<�(h��H+/
��{�վ�{�	"m�4)��bT =NE+����
qH�/��vo3��i��U�Y�u\�J�k,��u��-�>��%X6&M�v�]iySϔ���,M�;�M��*�8)�+�%���聮Ī:��P�b�5_բ��*+7VO�	z���������QQ44��.B�Z�U
��ԙ+[S�V����P��RHJ���MI�/R'^J-����q���bA�+�}�q����IHG&U�沫f�6���'g��ү�Ͷ�֭JdQ�~�G��p*����m�LԳ�ؙ���x�5���b����h��H��
8�^�Kܨ8i.Q��t���+b��物g%�Ju��۷G�tZ��6��+��)�rd��g2g,Sx��1����r����,c��,iї����jU�zr{��F|y7����\A�\�'�!SJ��<5 ����S�2H!��
���`�D.�x��Wd�Ʊ��L	��/o���eBdL!���;�p�x����s�,9��z���WFFt���֎Y��0�ڣ��$���������Fb�_��,�?�{T����v ��q�O3t(���G�d'��dIni���9(tl��l��W�����i�����N�H�G�1�f�CZD����iT��A�]�-cL[��JY������/M��$�l�:V��iؑ{������4-���_$XN�UN��^Ԥ)���_Ɓla?�O�ʊi�e"6 ]k�-Y�j�@N@$V.�?�{�r՟nӺ�(kU!�Ǫg�hA��8�{|���^��:�:0�ˏ��I=]��7�k�ӗ��o2�R���(��s$���Ɣ�Z�^-�4y���	i�2���=mh�*a��؂W� 8��Q����^���)S/꒔*-��ڬ��t�Eޮ���#\�S��*��1^�"<H���mm��ϗw1�f��ȴM����g��ћ��[X���X��L:�k2�JyY'�\Et���aX���]��s�ˌ�GHZ�(HS�?}̹D���)d��]T%�u�l�S������+~�w3���	����O;$�!V���Uɽ{9�W8+G6q�anlU;)���4@d;AF�$ɵ��rbk�D;'�;̕;\�F�2�pռ�Q�`Y�����,
�3�h��D@���eƉ���9m����a-��wy�9�V�ʷ1�O����m힄���is�����ͱ�%DHvg�z��-g 	��g���QhՎ�Lz�y�U���^��Ū����1�	q�N\��}�
\�n�����(����}���ݖs�%h�1�x���N>\�y@�O̿.�i�V\P���)Ÿ0gQ��G�"���ݑ9BL���p�x��:L9�I�JQ�I�����,V�
��>�	G�ն���'�٨��CV�Bvo���0��Ͱ0����W��q���\~��Wh�/h�S��Jw�@�kڰٿ(:<���h~r�f�Q�W��,�ʼ�`v���b0�m�Yq%����ԕ~�f������I�ò ��#��6��Fl9��dF��Ϥ���h�X�%s�BWqt<Hh���ʁD*� ��Uֻ�(�3��QT����_�	JF;
D�$��ϊ	>]����-��� D�2͈�絗�A����u�0F���YYYH Hĸtć�u�̾�?�P���:Za���L��I��@Y�x��R�"������zQ����ݒHɎB�������x����Os�6�X��ʯV������y�{h�CTro�yhK�C�{�N?Hk�^���t�3:fC�v���*��pAX/v"��:a0�>d��	���"p�pJ�d­R���{��ڿ��o�m���k���w�pm{�Hޕ/�x"9�f�nv"�"=$w�����)+�a�~��덋>W&gY�S����3��ܣ�b��5�;��� �77/A�B��Տ�#E����7��(�U�b�K��}%�(Y����Y�����_��l�6I2nC�<"�΀�D�i4!�b���~�R5?j��$n�Z���B^^���$�O׮����'K��Z���@<۽p�KQ(�y�v	�Xyup���6������7���t��f�A֛�v�]ʣ�o�:n��mP�=GwJ�?g�IR;���[7b�Z84�)���*H?�|�ne�A�?�U�?@���t���)+}�`�%�F��h�ɝD�ta�4B��ެ:~�&|�'<W�k�ȲWy�n;�'�|z��k�>n�����X�o}f�Ai�YCx![�`~�Jl8=DVO|X�_ڏ�y���܇C�%6N��z�dn����U�M��0S�XV8�@p	�)���dV	;�&�
�wҺ�V�ej�F-��P7��+��ߔ�-)˰�X����Φ�� ���O�@\��,v��:k|��.�8��C�(%G�K{�@i���rB���h�(Tۂ����fl͞��-�ã���+���B�3�9�������g����k��_�b<�}�op���0��[��,v�Y+����B�� �wq�"X��&;/H�'d��۱3�D���B����3j�a�_G��ѓ˷, 
�L>�{j�է�I7���$VX�����g��U?õpo!aP;�QU��`Ӷ�G8� �g��� �'�_��`9m	�g�>\�0�'�MJfY는��ŧx���r�Y �b�@�5��J��\�Qe.
��
G���(��UX��iu�(��ۗ�01�%��	~����4.bߩAƬ�M�׭+��XtgWF����U��c[Ne����f�`q*`���A�)el�tJ]���w�{Z���@�cD���r���hU�+��j�_�5���H�O<�ݬ���'lp&�ӼG�j�2ԙ��Kv=?��x}�W�x��0��o���+�Rɬ����̏ �)��9v���}���Nzr�.`-�h��;�ܔ� C���Qh��9��ĠO+�3
*&��EԌ]���T)n>��w��@q�B���9�)��g�,����AM0�q�)��s�}V����5��q��#�c{lC�J�z����铙EUZ�i}<ra�K1��������8I���`�����/j�n릊FF�h�����U뭯���|����s�J�����~��/�/����ѽ�|��i����o1�ں"�����9�Q��zaͿ\@tzsFSG�C�h�}�<�	�2� �Nz,X<4\��S2˙�8�,$G]69�p�z�e�<@�|�(Xm�pR�g��k��}0@1c���h
�i��#�n �(�Z ʈ��Y�����Rs\�@ mD��q�2 ���6������\_�ԁ��ќ�t:��Z�"R��(3���[&�a�凾��j�#u�N[�Ɲ�����v?����������5�+\��;�c�,���!�n�~Ђ����Ll%�r�f]+z�L%���eɜwc�!��J�r:UY]����(�Һ���H�B�m�n�������ܦ&��Lz�)d��/�:����5�M����cr٫dC�_��F*��T���ڨ+���$0������w�-hL���`�("V�����{-������5xa�{���zv�Q��{���ۯ�6�gۦ����r?�CP^U`�i��Mt��/�0-Aé.�YA�ҷ+l���T�o�Ė��j��"\�=�{�V��J�8Ԧ�t��>��fAd+*���m`�m\_�?�O�$zF��Q��2�ۆ��1ϲ{8^��5�����oZ�a�v�*>p"��jjK��7}��M�W?EX5Μ{Og��!l��&��L�Z����\�3=�����c'�[ʄ	;0�ɛ<S�������B*�d�N,\2ܕ�}�1z��&��K-�(jГvG���E}lؓ4��7�ۣ��������Ȼ�3��"�����?�����Q���L�s���.���u擰ӳ�J����e��0�%�j��A��i�4M��ˊK���8���ÖY_�%�*|���@�F���i���8�o
PU�i�s���Nѩ��2����-d�U���l����[,x�.�����f�[M-�R�9XK�2��ܑA���o��=�BfV�B���-	�G�������-�8��rO����6O�=��%u� F�M:��N��%�d�N��I�2lFHf�
��u:�h���|���Z�7I��	��3�a:A��UbY�;.�t�\&<Ċ���ט�=��-6�<���?,�]�E���̻e�!�|<-�,�	U�#vtw؋�}uz���z�Q :����%��x�m?���-퓖��R%���2*�Z-,q���U�z?�]��U�9�t�!��o���Gx��~������Z�5Q��S$J�?M�V�������e�Ψ�޺z�V�c�;bd��)����4�h�����BO�'���>h�/���u=��)��\w�j�G��Яq	�����˥�z���U·���	^鼌]��~Y
ʸ����zK���\���)e�����`���Z\uU�f3VzH�|��<Zd�_v���^Q�'P�)|��Ӽ �̛��cI�Z���(�O-�`Y���� ���]���z#��v�#�Ǚ�k�C�z�N���U�c>���0T*)�)���]e��'��[Sz�MP�F��1#�|}�\�$�~*�5�^?%�j^#�-e����0��de�B	�D�����Le�S�����
�-	�E��3��q+��x',����wEɊ�`6����^�̇��0Ay�h���[4� HG�nЉIe��\:~�}�h�5|V�9W/����������J� /n�C�B ����N��*AM�3�O���Ou&)�B�@t��E3.��0}��M��z��y3���	��U������+Ȧ�&�`�җ@�:�	��s��P�¢��u�g�Y���xN�X}�.¼A�*��|����4���1H`��"m�=����4˛)=���[Դ��-�>Ӆ�r3����dy��q,��?/�;%�_kF�i"z4J���ׇ@��-ꌠ�Xi�� �r��Nf���������g�$9e>�������'�\�P����ߝ�G6m��ڽ.閥
gŻ(��;���z�xi���������vĠ� X�CͲ��>'|�S���s��O|����FO�RGfC�{�6"�川��8�����J����H�#�>��2��U4>�dTM(�+���KZ%?|���O�/Vn�9�^�1ߺi��b^n��T�ٓ�?Q<�5t������3O>X"����c��#3��J\�*]f�3 4�1�����i�J�xz^�M����	�ZP��ʧ����A:���r�k`V\Q�ʲ�֌BIn���k+�5 ��N哄��@\}����9�7"���z�	��][!��1�������0Hw�,���<�;�Z��'L��g�Y���AO�4�h9��^�*�f��Q��rW�퀵襓!נga>ލ��������җ5��=�V���Wzw)�F���-Ȍ.R�|�`�����@B��]���ף��׳�"�\�m��������/V�FE��v�+(w����-<�Ӽ�!
IlV�����<c�Ra �1N�K��������v*�����Pq���<V���Kq{��t�P>�v����	�EKg$�̩#n����ؼ�h?z�M����"���ԁ۾H����� |�>���H�C%�d�qU��<5THB���
L�+*@ś@(���H��J��R�)���|5�3�D^"T��΁3��w��Uhc��:�=ś|~�6T+f^�I3�n{��ȓcm�p�PkdȘ�`��g�	��=���^Z�ڏ���t'�Mmq���s�� p։��x�O9����<����!)rcCz}�M\�����y����D|De'��Y�7�l���2�/�'aCs�̚^�'V��XC���:��5�q��cs+p/�WS�Gܠ,N$���ذ��"#���[��&C��Ý��WMD�.��5������Z*J��,�z��]%I�y���N2��8ƻ�V��V��S@�I����$��L�$6iT��O�6��ă��b���ل��û��b ��:ڽ��1)�錉ގN�:R�c�u��؎�c�c�B��4��iN��Ǧ������X�Em� �B�+��V{[��J��KŠ������\��`rq/�՝)������+�3  a��>�D$������߯N"�������7r�����c�K�P������K���U�0-���ATؒV�&C���=�FjQQ���,�� ʶ�ٔ/5���O�:Dz�R1�',esQ03:��XA��&@mT��d�;�ĭ�~��XwC-a�o	M��b�Y��x6n�#6�9��ҵ�@"%�1��W�3���m�;%7���::/ҙ�F\�8fe+l��S�f"�0��hZ|�Z h���C�ѳzJ��� �(���X�c��<?3�ONq�|.�\/��eC�ɏ�v�
�q{h�ۅS�>�B���ji~�#Qb��mn�-�X~22�I_Pb"���2�TA!k�c��%mk�T�X��V�l)��=��e�4]��w��@᮰�tr�h���`|h	hX<�ܔ�nA3����}�m��O�~��"�9׽$	[���8�����yxU_�>6O`�VJ��EoR
�@�`��A��k�D�^��� ����st���D��]��)=��E���O�W�w
t��B�2�D9��dj��|��~@�%��I5Q�+�l���u�{�?2=��0�h"$�̋5������JA�=�� ��@ ��#ˣ�����qAۣc#��ޢM���NVh�#�	���_�y�"�>���
_ʿ�aB�\�]J��%�X�rܘ�Eo��lj����EApҺXQ�Lkp�ۓi����Y���G�~����Z�9�+�G��<�c��i�-��h�E�%�����W�ǚ�� ��]�$�	yuY������Y{�"�0@�s�1�o���:��Ue��u�����V@bc�����Y�.An 40?��4�۩�~5֮M�qqVX�piNrn��}X[x������9�y�`�S�!�D��������B�^I�k���+�Ћh�2�`V��8�2K�f��g[���z�!��J@�q���������Ĭ��~[���n$��h���g��Y�n�d�| ���B��8-�u��pU�a9�Z@�޿�Q��<ig.?4�%����Ʋ?XT`�	�s��n�� ����v��R���U�;��>�~<�F�i�4b�����ݒ_#�{�Y�x��[2�����p�P�e�WG�p5E���G[Jzk��ʒ�}�I�J�����x_��;�Lڃ��[�f0Q:��;��+z��"-Oٴ76x\K~����Zb�7�jN�}�|��5��ީ6��r�᠊��w�f���`�q+ck�g�B@?�Pk�հ���x�eM��Uj��r_�_��~v������Sx��?�=���b�N��=�ʘ�h_�I��w��e <��'ӗL�W��A6�Nb��-�7w�2>"�%�����&ɊҴs�'�U�[���Nxo?������:SX�����,���ob�'_�=w�Oa0�����D��F�`]_�j�"�0�ѽw/<ـX��Kb��a�u��͎���R� �Oh�!L��a�{�4�t��C(Ή2,y0x#���Ҭ2[���(�CXp��?$��D	 &&U�k7@�OI�21DN��@=1��rE�%��:���st�|*�����7`{I��&^4NQ"^�Ξ�1~�<�q���[-�.���X�5ۧ�[{a�(���̈́�{1�N+I�ZWײ4��!86+F%}IOQ�����*�R��U_��R_,�oM����89)��:Bv����,FޣRS{'�x�m�����j�^���fw�z+�k<�����$n��/���������}�vg}<c}��ه����� ��M�c�|�4xP7��EᢝB����TҰ��C��wWy�����s��V��h.�夜�r~m�E8�y�e�CA"R�_uW�ID��w��|#g�L<��܏��U��ȕ�(o��_���y��i��R1�y.�1�� *>1J��/��©7����G��`��r,K�}�S0��G6�
[i�_Ԕ�P��w���+�S{�T���*���a;A�9���+����>�8f��~�_d�z��<tD��np�C��q�����B$�2A_���V*���y�s���P��UI�15ұ��e3��#�#\0�WY����)b��ɗ\���	��SJD��O�L>f��2@d�8�#��5���+Ϣ�k�x$����]�[T�ڄkM�7!ª�@ϊ�hڃv�]��������_.z$�6�9�c���'v�$_��S�1]n���q�����6�@��cm���� G/(HB��$Q��4v��KmuM��_1x�sx�j�2
�u�Gu��yVmϙC?S�QͲ���{
���W��k0o����@�"Sx���$uߠ�;4�e��q�f�� �d�{Ds���I5�,Ǎ���ᱶy�1=#�����S4r��[:4�*���5�p�ڃ��=]�/F�RqJ�ʘ���Bs�s"C��0қ����С4�EFm�'x�ܵ��E��O��l��j�����-8�gb?�u9�cKW�G�#�Os� ��s0> ښ��h9��̠\/����I0���ӊO�=#��'�!���W�v��wʯ�2�fU��'Bw���t ���eO��{������q�Om�o�md�5k�h�/����B%��ќ������t5^��L�q�������Un���z��8,⛠A i�ߔ�Xv£�r���xԚz�D�	�=	�u����b����Xz}��1��Z�WL��c��]>x�Z� Rk������{�!��zH
�ג浚��T�aB�}�.��2�[�,"�[�] Ƿ�7J`'�� ͷ�q���x����Z�H�ԝ�ҿ�`���<��)<�8�������Y 3߶6kL��V66��2��1Z{k�9�hRw���_%zqW�=�W-�0�	�2:�0������f��gњ@qE9�鬙�fO
In�6&]K#���V0�^��Ύ��}��՗	���Yb��4՞T���[�c�����p��p*�Ke�I ȒC�߫�4ۋ�S�[Y��r�\
l"jz'������1c�����>R�&⽓W�_�>�&�-��@z]h؛��"��A���&�-��1�����L�^쎼m7�>�1��uq�/\~���=o �$�(��h�q��:�ݫ}���CC�3���:����q��6�%�(�(�+�����(oz�Dޒ���`�]��B�����8{ zY�Ԅ����]��҆Z�)�m�}���,N�gކ�x�
	3�`7���T4U�1~����{yx�D9YB�^��/�A������R��]��ؒ Xx��!�JA����k0[勩-`�f������xmgvF��ڈ/Õ�\��0pEǏ;uh��un�P�R��!44�����L9�4��}����щ�u�����t�����r鞐Ζ�S)�����V!ZR�Y��������t��V�_}j����y(�+C(�i���US�PG)J����Ǳ��w@�ԹK��Jg��P��0����ltl���[�X��@<=�L"�e�+Թ��y`.�g�dkk&*����y�{���K:E��>�fͽe'��=�pƋ����(��_Rg��=�'��`��r���2��r�� d�|Z+�g!�[J�I�=�^��nH�
��M�n72T�DF+m��j�7H0Gy�DϨ�w�	8Qkd-���8���d�����5�`>�3C���`_��!�\^�6p��ɓ�L�^�B�ԥ��B���s1뚮9s�!�0�:�4��#�zC�O����w�K���9wQJE
�y.4��F�P���/(���rj
!s�xJz�̼"X�8y����?�x �� y<8�![T�� n� �(|u�w�cn��~y}e�R����#���+5�"���X����0�̯�.�{�6���r�,��!�%��(�2�>ԣ�+1q�	{��J3;�8�T�<����1q	~�yi$q�œ����0�d� ����܃��*�V��bm�2rJ��!�|�8��|/�.A����~��_�U���� �dU)��aU_)D�\�B�d_����>��89$FN���g�9c+�X�H5WEA�{,:׃�4��P둖	G�e	>�dB8�;�N�ƀ"E�~ݞ^��������n
e�:��� ��g��nRcQ{�)���r�������P�M�%��}L.jr����K9�'l,�P!�0�����4t;)҈�NtM5_]��i(�W˚���n�O�-F؈)#�����Ū��T��*���R�"�d˘�}-�m^m�����o��n0��8��$��u�>>rk�Br��9�J:�jƚ��E�V�F�͊� ]#!>P��,�d�0y�pU����;�:Q؋�j,=7��`��ە(�/�P`�mS`�ل��$ J��2��]�����W��Jՙ��X��2Ɲ�6�f�����i���rCJ��Al·'�KgB��eԆ� �e�35�����.QA�4?bJN�n�O�hG;=:8����
�j~�Jy4�d$P���������qn���d������q q,���]9Hv�X�e?D��9���c���@��;F�8.$ 7�G�����쪍�i&U۷'�w �G���`�xD�:��9�
p��t�q��i������#�%��;����imOGf4��]��rQ���/E�\����]ڥ�� ���CQ�Q���EA���t�N��M�����^ک�1����q�LŤ��c>�%'Y�~J�<G՝��YM�#����>3��p�����V���r�y���P����� ۰B����t�Y��8���i\V�r�$�L��_����(��.J4�g�H%���î�-SZ��	�+	�y���	�����Fm½��SE���;�O�3/yL�����A��8ܙMZ�	3�$T�M�N�-�H���:��[u�sT�0l��x�{s(���q� i�'L�㱡cܴ�><��鼒�/�``�ϒT軶V�t��n���I�ݗs����7�aI�̈́��N0�*f�T;g��/��9
���%)a�Y�%2g	1��m{�����nҎ��7<dR�&���?���?
��c��w��#$� �'[A��� #W�A�1j���vذ�v��3B*����'�ͦCԧ����������/6��`�{WMi+zJ�56k�'�S9'	�ۂ�7���M�E)7&��YzA��e�g.('���g����rFA������4�؜1��c�)G2��^KB�k:��M��Yz�P�#n�i')m��F��� �,HY�۶�ٺd=6�ˏϝ���v�h�dϻ��~#����ХBg�9���ƥdJ��0�ʤ�?tq�;�j9�Mf���o!!Γ/]Qͩs7{r)���˚��\k�eI�zW.VS�X��]Vj�}���z9����e�#W�Pew@H����f���e������cւ/%��yÝ-x���*%t�L6�WK�aD/�_G��^�[tL�Unޝϓm^FR{�@�wK�
,�r�ߩ�^�!T�B�C(d�pU�a:���b�:Q���̔�r�@8}�i�S6�T�M�Q��^��_�ûf.--�b2&�_sA9+_�����T"��\���K1YV4�>؅đV ���@�����*ΏqKS�M�!�>g�i��d!����N�ˣn� Gp�?���Xx[�O�M���Wz�?F�BO%/�L�FWUI������e}���:�]�)�V_�?e�w6�=��p����?'��U���0�w���@��s�;��b�#l��7��c�H����ڙ�}�5����GynŬ5�iA�u2L�,�P9~����;)m�o뤪@XЙ��ه���_�1r�Z����i2/���5,Fw��9؈ay�>W�΋�:C?�Ճ�!��##7���x��b���j:�P�����= ��Ȯ۫ǿ��G c���#Cܘ��������"��[�3�p�A�,��N+��]��-GkG��w��a���o�k��;e~�	�=��)T.1G򖅱�$�IaS��ɟ�ڸ|r�(�P�c�8��Y#�� ����H�;�_+��+K��F�_6Ӈ��[���eķMJ��!��.y���)b0[��I��]3`����=�(�ʌ�;�Q@�N�_�ؠSeeIA�9��u�6ȋ��&&�^�t��J����<IC#ej��1�ߘ#��h�l@��\Q���<�amb1LZ�w&��V�(�|K��=�G�Ӿb��ɺ̐rQz��2�(m[�m�� ��?���;|�`�����9no���*����i�0:-��t�T�w~�v3R���u�z8!��:t�ݵg�-C�,'�M��ߒS<���X��hp����� F�R  ���	���A��6��E�l�m��9���%�9U���,%�,�A�˸�\Hг[�i��s�@{��O�����ܯ�Q����0��%@�{#��{.�2�ڴ����+��$E�HCܨ�Ί��m`�Y�b���C���ۮ�MX	���f\�>�:���<��;�Z�]��<>�?�հֲ[od��Qw�>FG�k��E�)�O�����u#)��zbk�??.� (��p)��¶�����[�R��q��:�Ϝ�G���H �R�	F����������z�����f���F�tƥ�Qa,��Y�������̷ܐ�t��4��#Ƽ��#�p�R}Qtd���:��U6J��+�ݓ�v�^Ր��/؆��?�bL:��k�E�?R�=]�_"�4��)^4�Yg)QXR���.��Eo�7�<y���WN%�U��g^F����
F��[u�Ŋ���`��������%��Q������8(.��8�7�COgL��
��-��8\8cG���4s�#���Ў���+pT.�Ԏ������\"��Պ��v�i�\��6�@��)��S��W�z��K��څ{��5*2'���-�G����~.D���54%CM�Gm�q}�V}�k�# ���r:�5�v���*��y���62j�xr��<܌�3>����T�'_E�c>��k�o���F����w|�W
���E��֒>gv�s�!�x��T!�bK��b��~��Z@�~2��� Mw8���G� �Dޘ4
G��Kr���B�щ&`7W�Gh�J�Q���ز�؃�mj\A�o�xCw����a-Z�u�/�7����#5Q���W����iX��Bjr.�[ d�Uw$1���۔��kO~�t�A��poov��'XfUL͌����t����S�=�f�TQwi|$��M�+�%��dA��q��̿��(��яcW��d�3Fh��
��l�[�}��I�$�S$�ifn(qF����M��΁���j�de���d�>C�j9;f�W_۱0�!����)w����k�lKRO�Y�!�-����o�ùz�@�[B��+ɣ���\Zd�e&�(!z�,���[Y��t��,0�K�N�'���w;�Nk7^�8�b��U���T�+���G+�����Cz��� ����;O���"ʰ1*��
�1��G�ɩL���ٻ�em��Ǩ���Z�"ɹC��XuF^7�|49�
UA��H��Q3o1��ml��!���F?R<u9d�Auw��v�/�p���R'�a����u_𷸜0�w�/=m�}��d��^��W5�Hd��~�9=4�``�����J�-Y,��~�n�OL��3y��[���h�5��ĉB�e�Z 	��k���j��o qx�E����K�������w�ݚ.,y�U�x����F��`��켃#����q��*3{��\ZUǶ���G�P68@T|��O�O��
�߂L�L�����Ci�����1)oݷ;_|���@�P44�����ˁ��%��D��&	@�'��巘-tޜ4��Y�l�g������Z}�06׽��,3
�s�MB>�B��?v	nb�y�v�"vʫ�	C����V<7���Mp2��I�xbr2��a�ye,���T�z��=4JI��o�Gb����0{�vs�q��k�*���h�z$s�tQ�Ϥ
�ǖ���H:��r��Kx��m��罃P�L���A���e����1X�4!���wZ���u��*���ݮ�Uu�}����mI7V�G֨R͔X�q���z�C8����~��#*R��[��SZG�YI�PP/'���	g�ĺ� ?�G+�Y��.n~�H�Ҫ��h�_�H���.��{��S�Hָ����&���bщ���:!_�gF�
fE��o?�������@���c+�5�_�o�S��5����@�ؾ��5U���}��KL�/�K���] c�E���
���˩g1:�����ha߉���X�io���c�����~���˘�)�?�`���L�SΕ�ob"���>�����1�-1q6�j�O��}�[n5�eސQu�%���+�ۉ�௅L��̩Q,��]����QN��b��u5�l�"=nG�(~�x��[��Bί�w)|�(U�7	�i܊��夾9�)�p�	T^�5w�v�n�S�|��NO��N����Rd�.؄���`�G��k�����2�d���?�X49�9��뀸h�p������Db��cPiЅ�+L�z '#��Ǣ9�u��� S�ȯ>�R��|0��Gg��#6��3�y�4�2	j��NU,�S���{�����8ꖕ�,�ϱ� ��S2�c:�����Cw�1M����x~G}m�݉�_@jm�8Q�^��>��}�/-Ŕ��s	%���/�!��)+g���u����^��/{xg��.tJ��&�W���Tr6�KM�0������\��B�{g�F-����:�(۴����9aʼ��!ө��FѬ���$�vt4�����_�d4�5��>}����L�f��b0�M���E��t��v�z�lǙ��U3-��������m�ͮU�Z��YG�026���	�L�e��Y���%�t��j�k��w��o�(e��\.��7e@����6_H�P�{M4��;(��pG+�:9���Ɵy���.�A�������B��%3�!t�t�u�T���h�)8��utS���6����00�;��4^���I���7m�s���~Np��?o^�
�Z6�R��?u'���{�߉��ߎ:�g^�g��O8���)~���HVr�5�Cp����(<�Zz��*����"Z��ɫE-ָ�C�����ͮ߱u��%C��[ۈ���G�?�S��g��U��`F�f=�ɺy�mgh��i> kS=��ו�K���M룟��W����\T�W]��	�[iQ%b�p-�����\�9�����u�a^��-���m���m�c9�ʝ�����mE�u��Җ�`���a��˵PB0�4����]��{�/
��H)d��v�8��#�#���WW��|~�~��n�"NQ�V*Ẁ+ą�U��5ġ��.5���ȏ��7�:��dEԈ���]
�(���F娩�M$�V�,�C�4��BG&�x�庞�ƃ)p��7	c�}f��72<��O�K���i"��i�K(4�WH�QssH ���1w^����Ԩ���ʪ6��&>aBA���@�mS��;�:�`n�H���TƠ���n������V��ֶ�!�")RU.h�B΋�[<S* B�u�Pw�0=Z��ũ"��I�o����Am3�g;EM_��1�d�N8.��{a�qa��c���F=�2�/�u Q��}��uS�
ڑ�![��Km	O�3J��e�����K�+�|Ul�YS%��Pקx�Ҿ�/���� �(81Nv�7~)��|�� ��^�V��8[4Mi���퐾���h=�8#:��_��o��74�>+BE#�/u�n,'��l�"�-�ob��$�|ow�M�SQs���\��7�DѴ�}�9��?��wAq|���Y��̯���%ǧ�Ӱ�nB�#Ӈ�l~%P˰���������f����k��� <~	3�H,%Ū�/��?L���~�D6�������H������>�3�����7U�j���$���H��k��2��O�$�YY��.@��\�6�?׊�1�'v�VP��I�!r�[����\��G�iƧVl�	����wO:)ʰ���#�]�UjS�Nn��@u��hfC�����7n�����u.��5}�{XWp��oD��b]�|�D�e5����Q����Ӆ�+�|��-)�떭������C
�I��S��.�jz�r5��EQ�.�Z7�[��Ws��X$����!��A�H�����to�� KeEf�-F猴���i�j<*��c�xX'��N62��m�@ll��v������0��=�Jʵ�ؒ���4��e�B���U�NǝI,l.������"������p�/�u�0�TIX���7�	ә�/�w��S/W6�(b4�1W.��k	�_-���?��k}�}PE\_����jqKz1�������6ui����>�ĥ��B�~����%��q�P�Ֆ�����q̿��#<)���+d͔�+�F���)��F�����4�!!ͨ����� lV���^����u2�ڇ�FS����t�8g����'��8�񍶈�>�y4Q�����������R|��"$���JH�_��[Y�뇑r�����CA���9�}���x�yC����8jsJ0��g�����"�h�ǘ�XZ�Ј�8���%H����Œ���1��RN��վ_�qxv��[���R��)�0hϐn+��i_;�q;�2i�����E�n�'D��]���k��K"��G� 8ߖ�;{r�ʍ��Γ��1��
D���"#"�K�-2��M�c��j�s�*���Fק�>d�0�E�g]���xfj����p"�q��{�w��؍7h>+`�z���/�ᰮ"��R���J~�YgR��P�g���u�L��p�龽�u��@�I-�`���|��� �h(O�8��nK���c��Hz�xRL

>��L�%�Sɗ%�aH�|(���r�����a^�DOD��+0���I�щ����� �F�1*�����h�����⋿���r<�ҹ�����^LuY��x_d�2$��m�w���rUX���:���B�UFCa��H%��d2���t�-8N��s���7�׿�$yx�*AWg6�ɛ[�벃~~0��ɛ���Ri���F,D7�J����Z�yOlepb���"p"��Qt���K6�(�>�Պ��7Om�Kϊi`#,�ιx]�)��ע@lba���uq���C�p[�Y& ���*I�wFW��j#;rV�������F�ʂ@/�g]# ����2&��iru�G=],�|vY����L���.䕴i)����(j�8��\ԃ��-�����N�b����A���T�M8{�R��Tr�yU�\;f^�t������\��"z�51�s��p�PY��Kݮ�tEҩڟ#;��	'��m8�-	?� ��%��>��;I���:��6���VE ���4��2�~�*�y���䇑�����R�V�75�m�K�Z�%��{�mykô�yl�}S���bSyx�{������-l�h�Y .�E�Uܩ�M���J��92�`/b{+w�O���oJ�[�P5F{?���0	Q���H ��{�K	�P�,y�l#��L��,QФ7�iP9�?���d������ꐜA?�P�<�n��>E��o��T�hW�2��B�u�$�{O'!�]�"��0�ߕ�]y��Y�ru��'�r�@�BT��s�4/7&I��}�"���-�MIPa���<�Ӹ�]�T��(1�ߡ��S��g�#�c?��@k�	j*�����߾���g�[�����s���Oҵ�}똱�	(|+�i-'��5nd��ke�LMs��v�r��TQ^6~Z�*�����u+N/��B޼��.]z;�)�?��6�p����eOc*D �"���w�-��G{(:��VS�Eq=��|=�G��yC�K�^���[�@k��������+T��T
�$�_o�q�e���P�k{b�`�,@W1&��������.O�
���vS��=�%�[ ��h]��#/�v�#�O��О�;r���Ht�~�:H.�P�k����ړ�C0�S�����y�z�
9	�k�O�v��Ɯ�����l�q*yj�I\ul�0��vV�Q�xߩ���
ϥ�M�ؑ�+l7Q2G��B��hM�жV��e�׽�^&��k�?�6��i�}w�h���A�!�����8�6D�o\;�<3���:ӕ&�A�,	D�Y^#>�L)"����z�;O\�?ӈ����ojPL�RB �uyԢ��,A��?Ъ�lx2r-O�c&��x��3.�,5��a��y�:��z��VrN�&ꇡ��<4\{`�\�`T�t2'�����0�EP��}q����6���h���ʂ�V� |�� *Ξ���m��)����m�g��D��4�����h�o����y�&�[O嗈�D�0�`�[�l^#��I�/Ȃr	�U��dzw!U�_r�/:`�jC�Y�v� Џ����It;����q�j�K���Jj�Q�ģC.�M��19;����
({`�g��w��(����V�RzҚև�,n�ѝ��N2h����ۊ�HX��q�����)�i�/�*�ᅇ�����O��?ʏ�a��k��1Uy��'#��/B��ϔ���vJ�ۀ��ǀ��R;̠*��,�Xpq������t�t��5I�&D&1��g��i��lN������$k]z:h��)ޝZ U�[	[�ݓ������6.J�8�clK}ob�|:�_
��������{�	�z�TD*�����~m�-=�U�C�R�a�^�n��Y`����;-���yn���ˤ�z{���T���M��STKh`�E?Mz��|��f��%N�>f�Q@5X�t���c�㾇'^�X��E9��ɞA�E�s���޻@d^�/F�ڹ
�������opI��Qϻ�sZ�"��ii��s�l�f�~�Y��\r^�;Ѐ�$�����lh�d�y�4h�>C	��
�Q�ŧw�;�w;�sO��'~��!�I4bhNl'f	zt�����@���΄P1�>�{A��Cjp�K�
�ŝNÌ����R[� �zJA��y&�gnl����F�ǓРi��������s'�Q�~y��0�o^��W v�DY�b�?]�\��׾H���Ŋ�9_��6 ��=:<-�Q$LQ2�=�y�gIl$�!/Ue�'ϣT�K�	Q"�\q��>�P�����#��6��u���wڟbPSl��Oj)�#s��MǾ<�	GH����	k�2��`�SŠꈗ��z�L�aH���#�m���vx��i�K�����l��\�w{��˰��k?������
��<��K3/�3~�umߡb���k1{1D��o�w ���X,���'����ɜ�q'#Hy�m�/]_���?��HYS�J�����b-�c;,�̖ȻD�i,�Ղ�S�sPI�
����f#�����ƅ�&�j�+	^%B\�`��������Y`�ߪ/'�"�D�U�U���e��,���8�D�=��\����O
p��ʥP� A�`;���N���I��$F�5���r�n�?C:�̍f��Z�D����Z�^�'H�{�ߟ7���9gk�H� �sQ����_*Ѣ�zk��\��o�X>00�㿌�A1��"p<p��LT���!:]!*�L櫞h5ژ{���-V'�ŔHM9\����J�I���͉Mڢ	 .�����D��[�Z�6��We��l�����5ޯ��I1�+��$�� �YFR�髆!��D_�P��"p�	�0���XmL�jl^�<�G𭼶���?�yٙ�y�-ȅ�D��r:�l"����q�6�����]F����*�����V�Ŋ��z�~t�Sw.Ԡ�i��հ6`: �O�D1z	���]`�ʿ����e1]�i+��Yݞpa����L�]�v� E���W(���߫g�H����dSC�-�f*�2O�O�;��nDp�������pwW�n��~����C��x�(��щ�Uf�v�i��V	��{JfX��٠��z�9h���y��y1�V��k��{�Rl�gԽ_�\��S?Y��gC:�8'U���宋A9��E%�Sd�չ7�e��>}G�S���|�i�d�a'x��,���i��p�M�18+ @�җ�`��sj�#�M]$:��6�]b�j�)����;�ܴ)7�\I���g�-�d���Z.��؟�y���� ��j���A�ش5	.�`)>(��ɷڢS7x����<�K\������Nљ�U<�h�.��F�䐧���y� ݞ��R��wa�<��=i�x�4b�3շ�ί�?��1�N��=>�Y4�c�T�_u�x}�qX���\�,���gSq��X�*��'��'���bM���~�R�4�w��)y��%� ���N� ����Y�����P�ǜ���
)�p��'� �F�N�#�	�n��\����Pqoٜ����s�>�D��ҟ����]E?���ne���Z�u�;�>E��y�v{�ƪa��#���-|sm�?��KT!�e�m��y�28
���$�N�����ޞ�6�9�+c�<T�mId�����T.��N�_���@�����<���;c*ł�tx��R�!l���r0�9��R��vH��m�.��)�$H��8���53�D�`�*n\ֆ�T�����j~t��	
3o;ȶC��\���#��V���x��
1�m:���ʎ��T�dc��M9�j��Ly�X���*_��^E�"�~��x�7����i?oH+	���A��(Gc�;+l�@c��%���f~	Ԁ�i~<kY�e�!Z���h��m��G/������TN%k�yz�.��S�@�4�Cf���_����n�a�����VWueScq��~=���C�����?�A �=�1C4R���>�Nؖ���c�^k��w�����PԨ��I�f�&�,@	+�$;Z��N2O����m��S:��O���;N��X�&0�>xk�6 v�9��p�����l��ܾ��H�� =�HC�پ*h.�T�~9Q�>�-ں����~:D��]���`%(ac���wZ8u9�4AYb�b�pppS�.����W�^��1CE��]ޥ'�FE�jp��� ����X�[�}L<�P�W�8�.30�aeef�R����η��4�]ڪ^!�me��x������e��x6��%�<�/ �hy��W��'��w�_�#�(y�֒���*S�CkZ�#�U��µ J'�6$9?�E�i�b���߄�B� �#��B�U��(5�8m?ՁmJӾ(����{�]�"	[\�$��|Z�o�m���Ę;����\��)�q��XB���@�s�a��ߝ��L9��x���7�j� ǋ��T���!�9�6FUc?֌/�k�hb%�.�צ<깐��0�Ɲ"̋��� 8Y��\��Q����n��'���q+p����j*:?ҧ�9q[4�Sm��+zQo�>���|��>�K4+gvBK��{�c�8����0����=Q��e 0������'1�����*�y�/�� ���B\�V�������)�QAƑs��YK�4�yI*-.X��]E˘@>�
�{1���@��(tz�T�ͅ[�B&�hV�Ld��=�6k�`I�[l¯�_�@mx1J�3ϻgE��ߡhQ��t�#'�������j�	g�k=[�����(�'��ϛ� ,_�����9�O��4��Oǟn)K\�SƝvu��ZA{*�J�D21�e����䏳� �L��6�ϗAnn�~�������}�v�\�?	�-�u���ޠ�K=l&�����m�s�&��e�a��#��Mgml̚l�&�%`YO����"��{�3σ�O`�=m�A��9B�>�V$��n9�^��n������Y��,�ga�f�2�7I�n��`�<>�������a���F�rX�l@�c���}��w0}�"�J2?�L��3f=�?��f�z��4�6�S����ݫx����-1�~R_Ne�آ01����/~�x�0s�93O�"���Z)`"��\"�Ϣ����xՋ�:Z��+O�Wx��ޥX�  ��L`�|ZiS��]��9<���-�U�-�?�/�|a�U�0����Kiϐ��Hb܂h�V�} �����Ny�K"b������^H�qpU�gh`���U"%�/�}�9U9o{]Y�3&��j/����Ekv����왡���ǏJ6��R��cv���=����(	d�ڌf��]1� O$��x�#b�'�~��ъ�Ph�$s���ъv�a�g�W�$m��*Ԧ��<��^��0u�ǫ�y��p���S�G(���������9�\x�˯<�|���:m��r���7T��!^�{�u�����,���c����#�aS��&��]��=����#�^S��CN4h������[Ƭ����pZ��F��4f�������
_��>"/ ��^y9m�tj����إ��\shI*�z��m���[a�.��\�\ d��ҝY*n����� ���A�xB�G��2�\���TP>�]L&���>�
2�v�f����e�o��4E�T/ɝ��W��(��U5\*���w)@{��ۢT1b��Թh?^��h��YW�ɍ(M��m����2�ÃC����C���w�}1w��0�~4�p���Pm��d%���i��ʙ-�]��ǒ���5�3<b|�_S�0��x�7Eu/A�[���.����AY�8a�,H�w��~�MFw/��VX*��-Q���� >?��BJS��"����g���.�
�\|Z�h�d���AN*zw�P�l�{H����#@k_*V_��-
��J#_���{Y�^�v�������ƘkN�Z�y�ej�iX"��ҘxaD��#��{���<���ivjі�w�9}���֫��>!�rH���D�f�R[��կ�>=�ShP �{���M^�����N���e��i���۬�Fn���-�K x@�*v������+6�HO���)sv~�
��T�l���,SD�H���M����*����#}tWbΠF���p� v�h�x���
��+����P��C�"0!�a�G�^Q�T]�`�,�l~��\#�3L"ؙ�)�HT���{ �͸S�r6��`g�$�������?{/�z!b��̓��P��C�r�
a:��1DQ�Af��oH	�$�+2�Լ0���͜Lk�Zn�k���e�Xaf���Zir�Az���H�5�J��lz��u�s%>�fG��$([D�E�*�8h��O3ǁ��'ji���z��wZ��z!S%�����h�F̬ᄐ]^'�� ,�V���LT�$Qff���;�n��k�u:}>�y3�j�7��Ԟ�L-���%s�c��r_�p��\�Z�����`�Cq�������[�OUf��[�gKQm��%ҹ�3�Y�##v)���N�1%)0�^��̬dt-j�ᾧ]���/��O?��w�΄�뼗��*�.�1��V"��D�\^�H�Y������&�b�L]r�⪲�3���V m=K�/�EJF�!$%�FAu���X߮t�"兾�q��!������KJD�ș��/�{{�c켪��֟�{�7�0鶔��:2�}yu� b�f�-��Ą;�KBQ<(+�u�G��/f,��f�L�ρ8�Y�D����a&}�����xv㨬;�&ޝ얈	4��Ίr~� &����4L���ۮ��E��S�p��#sC�CR�y�维���P��"���~�c�X��L.b�Ę����m�����yH�K7�1�.J�6���E�fR0������'i�ŝ�%T;�iT�)��qR�4^�3
O�
�bl�k�����mK��z����9�������`	>v���Z��'�A�s�0g{��� I�цl�{���rf-"� ���;���@����-�I��7�!�uS�3S��JW,��Ԛc� <�=T<!��о3ҝ�f@�+Ѿ��M	qxʗ̫\r�z�?2tl:!������p��k�	�w�S�������)t�M
�]��˩k"A��=<?�;������g���S=JuM�W`@_�@;���0tP̡4N�mmN	,�ʝ�ĺ��dPp��EH(<&��� �W�`���i���зi��M�>6T)�)r�Ʋ�)����c�/QO��5��q�A���,�����M�5؅7a��[m��iz�ϻE��rH�;4!��׉��a�\tƺ��v��	�ݒ�;��2�߻��K ��x��`]���$ѝ8�;^|�����oAf�;��T�1�B-�<ӈ�"�\�0� �k��(��o*������I�L�(�Y��*�6.vh�<2
<���.H��1\�Fr![S�P�2VPf��L�'y�3BX��D
P���
�s��5���>��w���^1*g��	�6�x?�"�Fk�e4�E��Ɯ��T�֔��|`�.�OHL��j���ҲT����+
m��I��D�7<�hf����7��O��&u>bK$d�ξ-u�o���dw	��ٴN�@^M'��]���y=z#�?G���VBpy]��7-�dG0$/�	L��戠���i}u�Uyy�{�MH����6E��kĜq�>����j!�R`wkr?��9|tN����V�^᩟IdXg0���_</�� ��0@v
������{"I��*(�3�ǹ~�����^�oit�Uw!�U#�[,��̳����&IH�c`8o�� �Yf[^� �_p6[�&�R^k!��ϋ�ƅN(�El�KgRm��S���qƧ�)�qo�9Xv3�g��z�,\�ݳ4�f�	�V-�O��w �ˍ5Dh��Z�nx�r$O�;�7�FL�o�| ]���xW��]�%��m���|d�7}�lyQ�</\.̿U6{��C��\G�f����&����{BU�R�� �id*�hnO%�%̦��T�g���%�y���H�&C��7C6t��P�4z��H�dJ�Z�Q<�7�0���\^������S�d�nH6��]�-�Uɟ��#���L�^���։���哣�M�3���_�s�F�/��C �m���O�{����2̛�Ӛ}VB�$�k(�K�BL�P�,���!Q��:�~jw�*Y�#���F�ؼ!oQ����o�@!�����ːp��U���!��&��%��'��zN�Wm!�&����7M�G��Ǘ`h�[k�`� Zi��S����--yK%	yҷ�$0E���.7ٶ+#�F-/�dD?}���N�倒=0��g��~���O�e|�X����r|8'+���,2�m�%u�~�qw�x*臿���c���=0\�ܽ�rG���΋M�]U�CLuY��]P���꘸->4�E��b@��4��+ۋdX�.�U�h�]W�xT��yp�?�A���NϿV�"g�a:��4TJ�C�K�2�v0#<t���(�|�����i�8�Z��ro�V� 1DZ�,��9�-�#U#��r�8f�ur�W��m��nv���Eq�6��Z�UW�#T��4�\�(f$j�ꃷ��_�g�(h�om��9����B�#$�sKgdvמ)~����+F͔�J�؂4
Y�=TBe�5;'�n��Q��	i�OL��cy�>������W��s���������JJ��8Fߴ|5N(����&��n�Ŋ܍�ˠ�K��0k%�W��|�*q�ù�����z��%�'�a@�&�fv�9vǛ��{�)�Fq��d1���$%6�ɒ/�ǈ����A������ߊA�vف�.ϝJ
�������SQV�E4����"������5DA�p�ѭ�G�B{����.��5����,ߵpD8i&=��l5�/���mOu?���.b�t����
��I �qvn�7)���Q([J�����!�99��x�� ߴ������&��Ѹ�2�>�z��M���:aV =vB`�L�ѷ���P��!�&@H�4M��Czfi[�3G?�����g��	��f�Z�d�܈�k���������z�rͻ~�~7B˃������L�
�1���L�bX\�&���?3�n�M�PVݏ[���2R�̼�Ygm�5C1��x�D~������B�0�����#l�<�C�9>T:N&�{�j�l4|�n�1���'j�;K��`��\8ʯ����#<=k88o�-��e�$<�S׭���M]��zm�Cڔv���?I��A)���$������4���n�tc�P���H�O7����{�!AW��b��ĺ�4��P����c���B}f�U�q\#�ci�A�_eVAJ���i?�C�'�J����q�]K������o�� �U�,>LZ �n���1��A��Ο0��$��_Ӆ��t��s=�L!%�	�3f�5�w	��Ӌ,���r����I�X�	�����~+����� �o�C�Y
=�o�2��2ԤU4¬[s'�<A?��I��"�u��P�����XIݲ�w��u�t5�\�����҅-'�D���W�0�|{l^�w�]�-"��1�D��!�\����BA��U��%%dl?��(��)T�zBq�ǌ������֑�l� |��j�%�����+M�8.R��D[��@&^RӁ��[)K�*y7�=�e]��T8�۔ߝ�e��a�QL�"��j����D����?+R>�v��u���,�\������$�R�)�c8���qr_��f���PJ�4wg]u?��H��CY�Q�	��f<4��y���z-���p>?����������ĳ�O J���n֨�i��RE��7�9~�? a�P����T��P�L��^����2��X�EC������k3���R��=��_�<71<fY�I|��֋T����Y���*�(�,���Ɲ^��t�w�Ej1"m>�1��7A)bb�s�t� [Oҧ��&U�Ny8t��),ɤ���:�_^���E��`���H�$(Ա��鐹��'����� H3:����ˋ�	��Z��:-�F��+��6�h�,D:s^ByKSa�EIw��FFg�ʳKH�M]�>�Ctڑ�w̢��j%lb8]���5�i���<DD�N���\�ҳ'��C�3U�׻�9Ea~�D[�����X��m�aN���Q�ՙY���J�+	��o{sTD��?N�щ
�g��R�'�~�շ����?l�ʾ)�Q�[]��ò�Z�R���ơ{������y�.F���͠�a$R�S��3)��Ҏ����:t����Qm��yG�N��X�����D����n3�,;�mL��sV,��������J�2���A�X�x��*/2D���c�=����L��L��N��6S�i�l={��}�f����ܑY�/�y�z7�(c#i�.IK��I�$6�'u/Z�v�w/�3_�� ��"��_�0��$�S�Y�<�X=���?V	�ɗK9^�#1��ч����$yq��<��
�jXw^pD�7�e�My�1 �����>����*���2�_M���#~D��^�m�$h�'�>�%�ᓤ�h�!#HҪ^;���-H�b�0T;����u��P�ܮ���9�y�a:c$�o�?-�P��n[��)RJ�����U�k�0�/�����
�3PY�]�o�dgFN��8����J�Y�{"�\DMn�����H��YV<�儀�٩?y49#�NOT��z��|�?)�����9�K��'k�"�8
z��t����%�J*�)}�X�Ռ]Ӹ��	Y��Bja�L;���V[��D�̔ڤ���u�]�Ғ��"�h'k��U���.�A!u��m��6�"�Z�
�K#���˪��;B����E�@�nq�Aī�
_��Ǩ��I�8 ��XT���Y��q�Ϝ����gm�~�w���Z)΂�4ZӂK�>'&.��9�-�{eL�3(u�WڞF)��������t��� L��� }�w
s.*R��ﴠ9d9H� 6��s�\^h{���3q^}�_z���CA�VAR��'M�6���� ss'������B)p"���2�\�8{E �к�Ϥ������/-�����Y6�B�/�LЗ쯳QR�� �$7�̖S�S�R�}}�j��+�TrZ�VamXvT�	�^��6eX$%P��v��R�����u����� �����
c��u8��3C�1�����?v����$��	8���^�- 617�i�矿
�l~�t��k�2�K=~�Q�,~�ŀ�.��6�,�97kj�ϲoxd����ވ�p&8�!s�<:�Y�`�^ ��sfѴ��;|�+�\��{��$�&k�"��k�7�AFh���!W�ܸ���� }cO�0d�T�]J�ғƫ&M��$N7edQ?0�����׷�}Z�Q�1j��L�+��q�lG܈�NI�GI� �,���^�P����i�#��%>�� �f������D�5T���?�7q�}��ʍ�6	�cEB ��	�oP��k��V����
��Z�x��};��F��i`Q]��ߏ}o�$Q��$w��Җ:�B&x����[��R�X��Y�}�� ��v4K�6y�Z%p���p٩��iy3��ķ�+�nRa�T#q����Q��7��2��:=z&w(9��Lz��B��RD�N��?T�r��/�:�7,�oy�Gdt��sm��+2�°~4�jQ�J�p�4�����O�)��@u�o�n�a��\�VkD.z�$L�i�7E7�q�!�a�NB���;seO��K1oP�Y� �Ǘ����'���B-����c�8
�V{�2��$���ܲ����R#jek/Gw��v�{c���t�M��>=���M /�߸�G�f��ZY��e������
�6 =bBۉ�ܬ%��^Xz�W�|����~�E�7�e�[69�����i��@�%��ŸVʔk<sxv
T�iK��q��:�u"��?�-Lt�F�T�? �[��J����wo�_~�vA�4n\,? ����,$�h����^�A>Y�w��-�A��^̇�zuS����,�~n�xp��3�ΐ��� �n����&�>;�*rJN����x:��r5�ԕ�*[����ԇ�qZLFyu~-�J3���W���UWPL*@_)O4TA#e|�������Hs+��)d~v֚��z�����$�/���IGo��Y��#|����-�1+������e���.����V��ޭWрH��x8��d6dm�[eY|ud�H=(4%^ҷÅ�W$�GA�=�x���?�ϱޕS��s+ =q�i��Mi#a��2x�?�[0˝q���mU�ïe�+��M����]���K��mU�ά`Պ\Wߚ6,'����k��t�k����;@d=@����$�(�G	Go�`�7�>�㞉,
�7���9*?�Si_��R�C 	(��Y<��&���37;����evI�����E�V���;F�S�?��fט�ˋ}�gC�C�>(ہƷ��E�kU�Yz����P��l�(�!u*!}�%9�*�C��� D>����px���<�j�ɫ��RB��&�E�͓sMҥ��r~�:e�7�83P�e
#)>��)�^��9�Ԑ%�ET��_|Iy�պ�A����=��'�l��i���ч�WJ�����Q������ψm� -U�N�F��ȩE��|��v:y�P85�i��� ���t5��i�e$��Ռv����#d��-<�6�����8�$�T�s�i<��e&4w��>@�hm������"y_�&�]��8E�R�A֋�������.���X�]�y\B3{&��6&�C��0��F�?}��ƟH_e�ЬZ=��@���X?�{���]��u2VN��h�9��
��j�U�[�ϐo�i�}�v��"���(cRvv
�Ի(��,SN��
�њ����}$���m�����F�R�3�@�T[��7~�ۅLm-�EV!2"��z=։��~���~�X9�](���.��Y!nj�f(\���
Ϳ�1޴���`�:}m�I�U��L��f0�#`C���Eۤ��v+���Hu�Hm��oPT���yw�� F�)���YmDo��fY`� o/A;�2�o��3�ۜ%^����
��1R0.�~�d/Գ:��k���-�o�e��%�Nkxa�E�֖��q�B�y\��]����.���A^Ď��L�9�7}0Y~7}�X�S��
�.Uj������vv���;�P������\��j.���{��ق�<��-:O��|Ƀ�������
	Dك�j7��ȧ� �P��������f����1vzQ]cÏ�i�Fؚ�B�
���r�>&�(��zw�m�J�Q��Ve)8)�,�f���A�O�VW�w!�cHF� �� #O�(oG�i����!Q
R�.�ъ�	d��z8��U��Pv	��g�Ʒ���JKjQq�6��d$�ib�ll�2fF(?�fӢx����Q��(aȒ}�D�J`_�k�Æ�Y
Ү5�Tᛖk���8
O��\(��A��.F
"lA׬���E��^�m�daSB0,�?���[�w�Lu�'ȹ.�"�����VØy *�i;������|}������_)H���$��Wnu�&�$��e���S�]�-
\z.Ч"�TeQ�<�:,U��>�ԉ.� Yn,��7�pG���i�|[�٤{cTu�Nԯ��Dx��?8 +����3�[�G����>��}�����0h�G"'��mt~t�,�݁�+~.�k͵��x�qd�j�!�N��S�s��
���~1;�4�Y���5J�1Ok��3�)�S�n�q5�$4A����vk"�fv����V܌Grp Zk��_ �C0D!�Zl�c��`n?�M1��B2��i��(��j��ɺX�JRÆ{��}.�KuP�E�⧓�B֎��71;����.��w�=f�I��gY�:�fH��N���&�5�'f��Z��������
I�$|r�;|��U��Ͷ��\�6"C��0�d/��.A���, <��Is�sL���wC1��8�X��X���i�~���p����f����֋9�6xVNc#!��0/	�0ԟ�7�^�ڙ����<��AA��Ƿ�݇{簺x�A樗��]�h#���(����]�T�	�N��{u�9��ݮ���M�u��eq��(�����uf����ף���p�[Z�����&�s�&���s�?[���9�fu� }�Nme7}����(��>��� vP���iM|�<����bׁ���#���?pZ�4K|ț3�Ø,r2�.P��e,�tWv A?#��2w�QzVw6��3S[P_�nj���y8�����`���;�y��M�`1�A��D��Q��'��ǅ͏����S�+^/ �� 0)֛LEl� ��[��GrI�u�פ�ي��X�~w�b���T��'���.m�e�&jΕHQ�� ������
�/?L���- /R�x{P���s:q��*�,����͎���h���*�B^��ϳU�;]=��i§���z��$�e���=32~�-����8"h3��Q?��b�&6[2fD}/��l���Q*���SQ,Y���Vnm%@䐱�dW�0pA׼��ё�17�ưe�б�R}�4P#-��df0*QDb�:Bjh�$��e��S�m�ր�t2b2�=d��x4��o����%`�E��~~�����!q�R���F<0R�E�w�V���	�JN�c%��6�n��D6�k�f������
]�{}�~��=��9=t�������cu6,��:�2u��}��b}����{�$J|�;
I��]���L�-��F޸}YK�S#�M�_=��Վ�q(���G?� 45�oq�_��s`�k���E��B��e�eIŨ������Jj]���k[W)x��5K�j�ҍꇽH�q^/Go�g�+ҭ��/ΖRΓq�hɣ�����t�I��u�ޝ\�Obmb���(�{��n�������2�J�*�5�
�O�:�'J�����)��1�g�f?�5�࿫k-�dg8����)�axɸ��;��b��0���K���C�����+3h�J�ϺW�{=_
XЉ��q�jٹ_�i�U��Yo�c�W�� ..Z(j���x� r����m�:�>���4�K�������/P�p��������4ŵ'~�0�S�Lm��J�D�Mo��Ze4@�,6|NLuL?	�G̏D��޹A{�������.���*���KVF O�w�&l��"��j¬��֚�}��'��jl�Ks��CYr�H3�ڸ�yʻ����/r~�<��"��w��5�+�Rj�v��Yi��!_U|j�Eus/
0�J/�<'�sg���k�.��
��y+7��SQ�xÂF`�W���Y��G��p �d�1!��D�l$������N@vڛW����4逢����I��p��m�Ã!�~4U�~������T�J�X��.n���_T��i��y�[))�w�2���4�5�i]��w��<@���#�����	a���]��%�|P6����g1 �t�բ\��~V�0�p�v�
�o�W�/KM��3�lw;j%k�2�q����;Z�|Ćd@� ���� 4++}�{�=�\��H�.�i��	�Eݥ�w
���.B^6 \��K���� ��uքn&/הY������wǢ\Q���|;}R���=���6,�!��QŠ���p��N�(6@mD3D���_:�������5�W�����@��Y�I|�X��:�$��3��J,MD�x�q��;l����2Đ�́�th��V��EL����"��i�O�쪗8����:,A�B=GB݉'�@&���f��� ��u��Y�?�k��X�DDs�2�T�P�n� ��\��Y���S��7��|M�7}�sΉ��F�Q�Y�l?��w�]���Tj|��]ʙ��9&\"o��*~�����h��k[��-Z��T��PD�j���]���'GPg`]N�R�
H2��Cp5���+]�dZh!���+/���@A���s\�3���74����Gl���P�b���&����&Ă�����yA�ȳ1��n)V:�X��}��˽�i���eT�#qeJt�D��QX6�+�o��#h�l$��#��i�D�-��-�\e�#������Ǣ!�$������iQR]I�~l�Q�� �C���q���
>��x{U$�+�F��bn(����@'�����;�&}�rw�����Ax�G���t�/L����pwҭZ@���j[������_9_���晫)��a��v�x��R�"���S�7�F�Y�JD>�5Ws�S��7�~ ���§���a��e���#��T���
XV���4����z"7&G֡�*G*Ч_��D�޷��z]oDG�|�`��H;�����P �2��c~X��<��7r.���1һ蒶���}i�ΥG:��cj�	q���=(k���F�B��S�N�k�ȃV
��m70���Y0DP��<b������X��H���z5M�_�=��6�s�%�&�KI��7�AξD[f�b�K^�V��k���B������4ä&�9�)
D@���*���-�̡�3�i��!Q��j>]�"<�ԏ�t��a�	#�����H�N�ů�_61Dё/�]ըL{fј-\���u!�U��]�7��8�c�i��9�B3
�y[T�2�����?�����z#�[��Ň�L�.�X Gʠ��5ݛ�'����mˈ;�ӓ,�m�Zx�
}�&���S�����ڼn"vM���H��` ���1�����}=������C yv�r�\�E�)|��fl�,����{7]��!�O�gYY�8{+��:��V���)�t�%c�q52o4��������BA�4"��O����B�I�������Ek{�w��ŋ�)6P�	��zG�:uN�	�<,��f,���mӔ��~�&@�g�����g`��=�J��R60���PB�e���}��UD�����L��SuW�Q�j��b�G�{lm��\�!:��v_�&�y{O��x{Y �������wj�����B]6�1�g?��:��R(i��("�Ӭ���X�2��#�3Ԟ-x�;��`�U�nY�B��<ȣX)�c;�r�����3L�Q��~j��`�����3c�J/����DRUQ.�����rB�I���R�	]:X3�bv����!|&V@V#P�U���П���l��Y�C�e�]��]TƆ��W�A���֫i^�����
��0 ���b�Ǣx�o�5���$��r� y_�c���4�=�n�B�x�s�b'PȐj�
Y��V��(��讚��gl�F��֮��`M}=���&�L����Wt���3,�:���܉xT�b]-{Ø	;}����mF� b4���Y@���(�x3J�Q�R@Ҍ2�:<z�]|��k�ng���z��Uf����}8�?'X�o~l#c3n�o�R��8,KR|[�퓄�����K�ϤB�a�Km��ܥb��,?hKd�!.�� ��P�A�Ҳ�������Y�zV��J�o<7d+{3�/K\��H�ȱ�=Gb�h�5_�a<T�Ye%��UP�Əo��i�L��O�d�q�6�K7��Ko��%��_����+��kz�u�!�wp	�,����XJ���H���M��TOȧ�ʚ�A9W\��y3�
�$V8���A�o�7΅4I'D
���p�����d���(����=��xI��64�Si��r�����=�Z�h���,8��M���Sӥ�>�iM�)�q՟}�1z�'[0|.�孆e\��Q�����j�I�f��x��+�e*�<��0�OWm�xV�{�G$I�]1���r�2���Ha��y^;�ۋ� �m87x�Zf_H����Q�E��.o�`;���4���;���������pp���B�a
Y�rB�&��D@��i�q5,q狉���J�_4���C�<�?{��Pő��o�%9&˶K|��kx�:�-�9�H���A�ZJr�#�z/�Z�:��'�V6��'q�a�����
�Ǵd�r0��Ev�����60}I��ir�3r�WLF�AO��;?p1�z�����{�]@�ImB�M���p�3�.>Π�����\���.p�(ho�t�{O�����Nr0�J�VE2���qm��'q3�=>˿��$�ɣCF]Ɓ�F7�Q{���>�1��i��?�)���h�7#�x}��S%Y�a6,�K�ݶ��*xnZ::�D!���7��[�.śB�'TR�*	IZ5�a���m8ch��-5Ē���<�Du>�`|i�<��_�3A؁�R�Y��Ȋ��f p�J���S�D��
j�z�rςE~,Q�};@V<�u]m�b*��%'�$ټ>�(_h�R�������:�<9������oI�?Pj/%)��1� ~�HU�y�������G���4lM��$J�BF���05���m�����@	߃�#��)�W�w�1�rC��Q0��=v������tniFuѱ�K��<��8��v�Τ�!)��="}���l�Th��M�T/��/�-��p�/�Ta~���e%&���9�;��\}S@�Yۖ1?a%No����`\x��%�����a��SvQ������*m���&���Ȧ�O�TW Eמ_�շ�H�����/�g��͊�K�T.�>j��ܡtҤ_$%'���lγU�(иC�*�_l(�ħ䣂�ф�-sqIh�dX�C �Vṥq���)���u�hgn�4B��6��T�܀|眺�p���r�#�D}e�i&���l�k�4DA�_إ�>����=N��ty���S��S�[�U��M�D��Н^u��'~�n�t�c����ϣP��u�|���� �&��'g�X�$=���X�Y�:��M%�x�.T����l&I�I���?@\A
h�Yp��cK�=ыva� E\�#��50�ɣ����r��pV�Ϗ;�#b�/%`��7����-��2>)!���LX�3 ��L��;YU#ֹ�����=YSȹ@R@�<�h�{3��xF��-��2�)��^���0' {�]� �K๑�$����Ѱ���T:q�\]&�ѫ���q��䶟wA�ja���j��@7���ǜ�I-�u�=nfU��A�ꞧe����>*��1_���Ot���U'�T�e��"&�bW5>�rAG f 
�f��7F��-�*���3:n�r�=���Q`�/r����T!��ja�B�0�WY�����ZVӨ�PT8�l��>s9�wq$��1Tj:9f����	��'j�.y����P\
���'ft1Mn�G��W��.9I�9\�׏vP��
ȹ�a)��L&�ɴ�@7Uk�g#�I�&�=xC9�by�[�u6x(IkX�����7�L�٤��T?� ��*&a��?�s�O��5��ɷ�l=f�w���;d�V��u�L�1�������[���ȣ�5S�A�mA��<��ڬ�en��Ҏ��+s���B1ᅳ��GGw�̐R�pL����d��D(�o� M�8f�oړ�b���Iel1��S[�SD�����F�:��4��:�R���	U�݈�`Ίn�A��>A��������˪H(P�������䮏ih��DÝ�b>i�JY'�VY��x=U�zR��zK��#����A�Z
�j��?����tB=��/���NR "���0�Ss�:a�2��W�WZ�]�)���6|/����3�Y��x��Z�<)9	�Ƥ/oA���.��3��m�Aܿ�f>>;ȗB�Z��g�ׁ�����iB�v=z5����]���`ϙ͓n;ptR���w��9H�o�nW�IkM�.�?���A��s��_����Nj����8�(�ڝ)�?�7����}�Xj,�*/����b��k�?D�v��*n����l���4�-�:�BU�p�� ��Ӿk�͵)��H|S�L�Z�Qm񶀹ZB�Vj,A{�?,�yi� }{�}�	sS7t�_BQ���B�Tk�fou�q�����Q���1�A� �_�gU//�b ��{!�)�ZN�����6Aܕ7H�
�j���79�בm�����H��N}p����~=	MG�jV`UY�U���𝤕�\O1^�4d*vXF1�]���>�:��CJCFL$�\��@z諧)�#�&�{R@?i��:�"�+��L[]�-VǣÀMK����GL�"!���㰉��&�K��e�C�2 �^��1WD��n�m�9����x���^����Bs�+������������W���Y�ֻb�_E�Gf�\0h4��F��#;i��?cV������o��O���Q�/�T�S�Q̏���M�T���	=T.=���\Ԕ�:=_�O�i��Y%�1���҂�B��p�b��
�R^���U��c:,�y �Ru-	x��48L��TO�q(æTW�)� �����%���T_Ʊڱ�$������Ҿ'ql��0c�����ؔr�6a�A��p�%�1�{�'�|*G}Q�Wt����N�?b�:��{j`��v��gD.�)�;`�k¿�v6�5���Xk2Z���/upEsX�V� }��W)%ԏ��g���pĞh�V���ܸް!ɸ�pRHs;s_��Y�y��D�������xRp�_�PE�X�IY��J��RK��H��R9���)�춼��G|�x^����y����x����z��g�l,A\���s�pv⏛-)��߭�~"��Dx�JPk��\r��*}�
޲Z����$���|�r���l*��SB�/��|:a[c��(Ƥ�N�Ulm���R�����`;��[��1j{LϨR�s��Gy-sr��MjG�,�,V���������8�ڃ�k��5�p�>t�iQ�)���ӭ\2����C@��gR(���+l��(�E����F�K�zJ�
W$��)��Lyůه^	�=K֥�sĪG�u�W��U�~�@ZO��/�Q�/��0θr.�ĥ��B՜�J=	@�ʇ��8�e�e�.���Ꙅ��P���e��3_�-.�B��tz��n[�w�@�؇+p��k�@��r���?����
,}���l�m&�r<��Y���Z�`�F��y?��5$A?��9�)y��N-�s@)�����7]t/w�0x7�Qh������tJ��8ך����0��<`cK����+2���w���%6G�h��p�X#T���j`��Z����;|��+�:�$f����R��PBi9 ��kv作�"�,"]1�z�	�?�I����x������wD��&�|{Q&a�I�<��Bj|(���!�_S�a����b��=hI�@97D�fz�'�����Y8iP����Li�p�4�m��A�*��&�.�o+����}6�c�^�7��.�/�o��+ro��P:!L1�b�v2��S�蝑l�k~���m�6K��ۥ71A���h��׳�1������XQ6�%�U��Ǭ�&��*.�d�(h`�>l�.��[�$$�>rЦ��\?��|���	�j����l�He�%���ҿd�2�|>�
]sj�1��P.�<�l~�ˀ��b�|[	;�;_lK�4���p�1�_���v���t� �)2�:�:�u]3T������Հsl�����`���$z�*����a&��Qӈ+`�Ka< ���	X�pq�n=�g��V� �h�2�㟭5l��2��4�B��Ȁ�HB:Ȱ�d2������5/�_��l�)Y&�;d�O3��|ΎT����&x����:o{�
1�n��Kd���lBk����8y��d\�a.َB�-�5����W.�8+K�jRy��ޱMk��sr��:�A�7%��Qc��U���Α�1<�?Kw���1�ǃ�]�6?{9۵'�r���w�oXu;:T\F{��6����±4fU��X�;�@�Y��y� �:3c��:%�VQn��)�4i��Mu/@tr�{iM`�j>�(�h�"��W#���da�)OR�s��!&���$�5^xn��XQʴhP�EMNS��K��Z���F��c"y�A�J��W����/��*�~K��W�iw��.������GVpʪ~�5}t]غ%0犌�W��+��㟜6R�*;�b��w�Y@kt���I铳& ��K��	��|~�S��^��j!I_��P�RX��̸�J�j�	2\�=\mZߔ>�՛�eq%��Y
�\tƆ�f|z!���1e_��I"ڜ�y
_���VhC�Dƚ2�<f�m��A���{-�����2��zy	8=(��	�eK�u���r����R�_
0=K��n�������=�#q��T�����c�WV+(l��l�I��7%3Z'��",�������wI�Ew��.8Tr�k&�E�iRT=��y�w��}�QCg��	�`]�(��.��8����C�˱A]	P�#;��¾uk8;Y����Y�6k�R�����Pⶽ��u���ȋ:q]&���Ą�x����c�.�i�6�]я7墷��.Z�\6���2h�����qY
GE�[��YwFX��j=�^f��#���!�0�{]�Kf����~Mʤ��4�'����je���H-�@��5�G�<ž����x���g��5�i��6��Dp~-���o� ���e� ��x�{��t�_���Ҽ�n�H� �]�C��>�˳��&��R���h��qy/��8���M��͚��'��pR}��|��5mX��+�_!��9�=��~�}��퇘�,-\������r�6C<D�����߇a��C���f�S�����66p,�|.��)[���G���ԑ�4WT��I
�]��9@T�@���4���U�����.��ɾ2���Ő�G�Em�Dc�_$)%����6����Y���
�1���qŮCKç���e���?���G*M ����wժ�q�O��۹:P {�O
	f+�d���|��j�?��֎�(��H���j�gu�(�q߰��\��g ,+Y��3+Fvd�I��J>�Mj�����R�{-K4�w��Ĩ�d�8b��4���K��
�.�i��U����u ���,'�NO3$���UԳ�x]X�0G��1�ćbQF�̉��(��'�{�.��u(i�|X-?�R9BM�[����V��K����� \��~��$��x@�%wu7M��G�hr��`��cnM�LP�5�[:��y�%�އ6���>6e(�~�O��bB /���y~��Wl�y'��S�9�����t�F����\i����@����}W(&�2��酋�(�:��=�숏\��M���q�!2�֮��ds,�{�K���k�Ķ,��*��ʁ���#��~�KU	^.����*@�.�!�Yy .1c2[s0q=��uܧ/�?y���� {�����{F����2ަl��σ{�>�og�ap*�G�!����b�p\$d�}���6��y��\6���J�ό��Sள�W�V����� �����
���ٻOWe=�ɦ��(�5��0X�0P�ڄ�4ڑ�"L��U^~;3��w�������תW�_�U����%ik��e����+rJ&�*��4�UW�LT߼M���޹�۟���������iKn�#X���R]ra�R��4��6�	�f�#�V/�1�$OF)S�b�)����1�)C� +���Z+�Z�f��ks�
a�ɌB��e@,ŧ�mi4E<��rCV_�֔�{�,y����gLX3o�
�H�y��:�f�џ�7�ZtV1�@��Tɦ57�hR殈�A���O��FV�Y���`IKޑ�k�gI�U�rs$`X=ǩ�?t���w	���A(���1�4y�����S�JNΛrە�2Y�V�C��w�ɇ��ޱ���^�p��o����Im9���������q5%9mkТT����עCC<qN���^�-��`���x���P�u��ɩ�"�Nt�� _��a��S���A�3��Va�#Am�!+�{B�uZf���{<�
��Yp(%�O �\�e�	�Ǎ�混��5:6���mQx+��j��x���Z��r#���,z9�:����Gw6v���fH3�)%�}��T ȑ&���&�i�i�1F�P	��1���^#,@�܇*���ן/���x�	�[=	����L�~������\
6�1B��ή1��.�bK�#mIP褀[�Ʊ���	��y*�6y �t��[�L�"8<�EBG�D��;��^�B�!>VP��=���~�$�>z����7�4�3�;��+0�p�殰��Y;�#��(�-��r��]�*bg�=$��?�ˣmSS��c���O�5M��&Z�����_ޙC>E��y��.�����  �*�����P���JJ5��^�� �����/��4�uܟ��%~�`[��q�&G�*
�����fr����0_#���0.���K�_�VD_z ;���0����ٵ�i+�x9�ial4��X[��r	qs2K�h�*��R���kn���"���,6X���$��_������_axw�\מt{����Md�J���`�p�������@�{-Tb8��1d%�>,�f�#t���6�#�����{Ѷ3��KU,O�.	�Ťn�$�����Rꚶ(�B��JxT/%�0x����z^�V)�//YBٗ��DM`�s~��+D�e�4���� �9L�Mɍ,�u�F�B� p暻O�]Z+�P^����gٳ��?M�+�(bB���9��̶��~��D�*[c¶��{zw�_��S#y�����_Ȕ���*P��Sq��0�O� �9��)_Q�$�����+�X�k���>iC�`�`����T���z�|v��I���3❞��qZ���R����9��\\����琜��!�y���,�yA���,v5��̜[��ٺ���0�>6c�X���C�`��nAz���z�@�m^�{a��5��w���B�#	!]���h�ޝf!e�.%�l����޳�2�0�L�ǩ�r��`�T��w�˽�T��p���E��M'Wn��@1��*Xt+�H4�a0���˝k%wF
LS���N�u�J�G���2(�m#}��2����ț�A��/���[�n����\�Y2�4������<M�\�9w(���/���pI�]��2Wm1��q��vs�aȅ6�">������OUD3N�o��iU�1��_0����h����_T1�>Rڇ,|��9�����"�7?`Q�� ���|����Q��|͖�;��o�Yr�!C�|-�(��0b�~�S2�_)cu7�j&��Y러�?�,0ȼ��1�vs9���	��t����&�(!5çn��(_�3/��N�X��� r�A ���g��A��N0�9�h��c����;����S�"2�ɰCZ(gk���r6����jDy?}� ���f�%��ţFx��	|���Ú'H���0�_�(���/��F��JK���~�f�����H=�\ѯ�>��4��%�$�l��J��jI:�"�Y��� K��986��=�NGM��G��/X���9D�c���*1�l?3K��Ig�$�벸�*�A�`��t�_��Ibn��JeQ��&}�%X���X���DD&g�
3�l	�.��u���[�)N�m.�P[�C��0��VDk��Vk�j�qj��Z�{Ϸ0�3͗�r�Dk���Z눏Y��~���
)���O�kb&U� !L_���ŷ�c6�2X�D>�����Q��\,n�X�Q�»ғ�a�k$�u�]�!��c��u#���w�j�27���xc;�n��Og��Hr�#��C�?U:�76W^��=���p� ~��n0��G�*с3|bد�
�䃃+E�6����!�+�!z>����St{�4��T��xb��~
���NH_�����	W3OdDzGcMn�l��z��rdJ��D��Ê���r0�:�|9�Y�(\ھǤ�?�G5�������{�ɘ�#_4�m=�j�Ƿ��'�IKi^�D�+j�!���l=�	2�o�R��?���ߒ$���5�)�?�o_��ߤH�>����S^�k	� �f�&{�M'���b�./-��r�^��z�f�}�B���31a�g��"�.{�F֚��ax.!�U��E�Y6�a��v�|��RS� �mv���a�d�ơx��qU�>�xo�`wD �J}x�i�S�}z�"f&����[�d���}�o��Y�:5�.oj�����e����J|B�W�o;��s$�&"�S��!��y! � �[���ݷc����d�I��G�H�nyӺSu�0(f��#oA���8n�����D��% U{�Z�5��j BV��?[� \�C(q��H��� �~�q�9�$�`��*�k� ��YҞ����yӿ�e�	0cЦ��D����#�ZүMa�K0�xN;|�ĵ�#�g(��a#��?�D�ss}�s���=��K-n�q�kt��UPZ��W�o2��@/���4+Ҿ�_[��F�0rը&�*}�׆~��/�U9�̚��-��>/mc�1�W=�u� ��Q�1�Q�M�/pC���k���ʝ�����R@T����|�F&&`V�M��P��{d��Lj���e)���{�N@?���*�B�2&��Qs9/��}4��`�޺/_��
�#XϦ��R$�ñ�Fl��6@����R�5����<.B˪sG�=�m����k���*�W./�9w)O=���M2���'($��R�5^�y�1�ס���l��t5w��6��Uo	!6�y����;�=��mX����2IKҍ��E��ު^q\�p	PWS�+�5h�����=z�ʲ":��nk9�!_��$ЎZ�1��~���������I�2J�h�ŶD��UX��{\.�Qr&��_��?�N`$\#���)'	ل �.��x
v)�=��Z׊0�ߛ5��U;�fV�gw����F�)F ���|RSa�&�H���2���b�ΰ���h��u>��Yԃ��:���i�#\�-��D�����ֵ}���Ncv���2�@��m#��!$� Y�\�y�K�tm[�ڽ�7/��6n�8��4Ϯ�'{�mP�sPJ���ڭ��-S����k R`�JO���~~:�838���v��-dW���,Yn�Aw��8>�8gR��sGYXNH�|�eפ���zcop3�b�OK�O�t��� C�|=�l^c[
��y�x�[�bB�:��ܑ5����`�5U�O�@��.����d�R]��p,!N2h^k�}#�b������>�VU�w������C��_$�]YQ-̉yB�����/V��g��X)�͌G$��!e/�8P�B|f�yu � ��t,�	N#j5^�W�hX(ȸ
}TQ����󟿝�&/-Eȫ�z�o����vrbR�)�W`G�R���1������超|-g�.�u}Pm���3���ӗ�AšH:�-��l�HrH����2I:<��Mw������{2�_Ie�ֆE��� �@�-�f�f8}�H�e@�y7.F�Hh%�1mm�g��;�`�[Ҫ}_E�w��*���C���Jx�����R�GX�6����Y��'��R��/>�nG]��6>�&\���ɨ�IIUI�������}��6�P%�=�OD�\�� ��5G��={�=1 lȷ�j��G�����Wv�z�[����)Z��P��_MPBv�&�W#DT�?i1�As<��v�Q^�	����f�w�O���7��Uc�mm5 ���^�]�Y���:�?t����ف�*pI��3^�a���쀶4�[@�O�­H\tع���:����[�>{������J����	mT��a��n��	����}�6��Zz5��`X��s�Mʱ!U�9Dw��#=J!di"���)��6�r�$[���R�jz��㋓�����w;Ԍ� 9�`՜F/IG�Yń.��~>+�g�0*��Y�?���U�f~tW�$�ீ�����T8ƚ4N7.��jp�%�7T�@
@O#c��m.�����''�U�4̮ղ�ê7�ݒ��ymD�!
Ů$S���E�?v#�40�&�p�6�{�W�|Dj��n��˓�����lQ�O5Җ���oo�����Q��Ց����ة�R�|�zm$��Xɢ2˙����ӵOs�ݷ���q�F!����X>�������?槨�˾X�'<[��a����Ih��Z�qx�{�0�����4��q�(����=A����_k�Â,R��[,&�b MgF�LWՑ�xC��n]���Ph�ـ/Z$�d|�ma�̼���B��sQ�6D�'�!�G*h�k���Nt�*H�����A-�"��NǍ��0��U������Q���/6�^k��K~�ѹ�����~YTN��/�7b}�F���p_o��]�yx}WC|�����xTQf0��W،ǁ�}`K}���k��+S��n`j�B5������&%:�U��v'��nϖ��43�9;x�w���f�1�uX��ٗEc��S�Q�-��=H���a�'C ���"�V9�D�kr@�E��@�{�^{9s��%E���ί�< t��m�DH�������8�Q+���,�7F�b��v���&�6*��&:s7��݁�T���KN�&���ᗣ�k��<���q�i(ϴ׮P�l��1Vv� �z7���N����)F^��seK�����箩`�֌h���6A������T�[��ŀ�5|����u��D�$W�j��Cd�H��vC�N& $F��>��RO2ܗ��B5�=u�^)���@j�#\�LC����t�ȳC[��bXt�*��X�[!my�K�j{�,����/ԃ~C����3�}]�6���Y-����GF��EE�8� ��qJ�7U	h9g�g��4ξypr�ʱ���[��fJ¨�l'�ϝM_��Q�]@�ą��X����w�lک�g�U4���G�� \�m��+,�u���vp���� v��t�Ǻh���2�U����Alm�hh�J%��n���ٽ%�8pk,m Y��h�b.�y���5Z8�w}"4۵��QA�Je-����'`-6U2[���Z0m��ĽX=��H��c?�� ��٢��ދXx�EL�V�NRG}�!վ�~:�"�Q![��åģHEĘg�Fp�L�A ;��W����p
B���d�g�)�yBР����c!ݩ=_�I����Stz-wX�jV�����3ޱ}y���3k]����:�j���^xe| @˴��zN"���Y@�X��J�r��d+7(�K�&����Z�SH��>�>�P�*�44��ޭ����I'�%"o>��/���e��{��*�U��j�"��f{Ǳs�����,_\"�����'B�%V`F���whR���P�_hUT�t�y�/lI��)X҅U�/�8���$s��>�=��Ł�p��9k2�-�������J�h`L~b|i���6��",�,c(�@2���b�������1�q��Zq����+����ѧ�]�!�䓘���=��,����K\�sm�Jt��'��B$��
�L�5LVIR�;�����˅�s�l�[�,G�����@T&�i[�� ��B�'�U=��Ng�� �����r�h������
�ryy\N�edcU�!Q��'�1�M#�=�V��	-�p���b-����$��q����$,���;���+�3I���N�U��mAb:tR0eN�h3���=��$��m{���
�J�y9rQ ����Bd�Ձ�1�qX�w��j"����Ck�������^ i�N1M��TFi0��c:���oG�pS�J��e��V�`
�_4�ב�`\�:NZ�azP΃U�p�������0�T�uB� �m��2�S�Ⳗ
��Х7C�z�h[s{p&���$׎�z�Oz�9�UI�S�0\���,9]��J���_P�V v�+ջ�_�\L۫T:[�f���l�9%���)30d���W.&@�.��#-�n��%2��'��:��nM�̿�$U�Ϧ�D��^G�|��4���8���ZA���"e��_F����-�
b�ǟ�v���@��v�_��Y�`;R�hX�(�-���_9&�?}���S�_��N�:�n��
��q�a
��Ӌ={FHsQ��S���*��	M��VjF.yZ����R�& g��X3��D���d��S�l��`M�X2�]�]o�Uf�����<5�o�y̧��!��V�z"��"�1�+��0,�����4Z�d��;
�k��G�'�)=��:���r����n�1uS'��F�o�+�V$"<Y���7r&���b�3
^�t��M;u�80\l#���
`���l�����l�A�Y�tl 1��d��������pY9ɴ�(n��d���x�u�鶏!"\������w�ǘ���$�XD�R�@ܑ�g]]/.����-���'�.!>ƥ��a�y��y��@b�T��O�`�tjS�Y3�P[�������m��s�&��f��YrɤW˶=���fs� \�B��d[Y���@�J�r��|`|��	�������b%�%MiI._=���U�m"U�{]�N �4G���`*M���7�re&�?��E���C_]���
���X��K3X,����Sb�{�6:�V�'�"x�C�?Xў��s>�\jV����R&�f�F��b���H��W��Y�ˊjo��0�aJ<�1�9?�������$��@��0yuCE�H��ڽ��\�0�6��Nl�/��D7�ͦϺ>�3�JO��� 
x��C��B���CQ�Mco�q���F���V;b�A�	��d�H.����f� �lT��̮/\��oA�ue�Er�e�'6[9�9]�ws<*�'T���7���$a�Q�JJ���>�a�z2@���>�qp�ǬbQ:��4`X.�{�Nlp�c��+����M&�D�:[�&�v-6[.���"�/�z��/�=r8��~ieZ����o9��
F	_/>
Z0�q+Zb
�`��C��]Wa,���'�gj8V3����Ū����k(�>;Mir~!��TC�?��|H]͹xˏA��M)�"FKW`#��|N$��F�I�����ڎ�pjꅧz[�_F� �p��F��a���y��,�_E��[��(R��Ź�} k睎�r�<u����o��N����?o�6�L&�9� E�h$z`�4��Bo����t�û��a!M;J �#�V?���l�n�
�a�[�������̭�L�fC����E������Pn��.�����O��5K��F�ȥ�:�8���el�a"�YKj*��U�l�Z��Z ���`(���RW�y��>���\:�q���`V�&��Ym�ox�9˸<H��)�\#,a���KK-��p,;��ls��ty��ua�S+��3�^��>�-(1%�o�˾��Q�䰃��(U�s��^]�7��Uח�
r44=�he!;@2=~m#MN�3�25�J"���9�!��#\Թ��qf�d���]"�7҅s>�f���M�P��\3_���U��~TC?u���U����nob.�{5��	L҅#!]�����[21�uF6�~<؈���ִ�A������C�����be�PMۮ����B��Z��9�-�
R���PW�C��h�� �*�.�Cl�@�j���#׻5�%g�P��W�2�����$l�m'Aз�Á��?����q��1�.^���7�a˟dD#��IN*BE�S�ލMѢ}�)��Y���"K�6�a`c���5��B[A36��Q���!$���KP@6E�	���`������N�eH*$�,��߉��)�p� ?.�ÎS�A�5�ȆW��"S���/.؂���nϱi��n�Q��w����l�)�kǮ�QpV9��t���h~<jCo�kbi���JI{|c���
��gl�q�OaU����Zտ�-�J��\i$k3Y�@��� �	�*��d4��2��ճ�RL9���6í����ߤ���=��}z@j<}���c�T��x?̈́!�~���>���TOi���խ���1�h>�o����	���#쟂��J,Φ	�㹦m�y)��$-O��!5��1����{�\�D�~\K��kl�$^-���޹�#���Z�}��eҧ�k(�9��D>����Z%UkJ�3�hjj�����7=�r�>�ј��`@'�Wns8f �	冉lһKN 3m�a�gDDi�]Hv�}�V��ps��]����Yr�>&�}�N ��Q�Ў����𶷆�D
�,/����r>t�>�T�%��*�Ubؐ�fe�*2f]�A���]��7�a��;�Y�t %�%�mR�'����%�����V�*�x3���^-e���|�t�c�Ȼ�ݓ�;y��!r�Z�]l�+|vO2.�2�D�D?�Tr��3O�{Ŝ�����VX�����(�B��8��}�s��ܵ��P�/	>g�89
o���+�K�~fx�b�y��'Tp��'r{�]��KZ�^^���6rO�Q����ό������N�������Y��ԁ��e%[����4��7�����薭;jxd��ݹJG��;7��\B��\����>F�i���̤Q�K����Y1=�C�Ȥ��n�o����D���`(O��"b#���2��-U�'��z/mɋ[��ً.�uGbU���OP�,D�d�_�pƱ$;>kR��Zu
-�f�g��1������i �:�����H����
Ҟ��܃���}������F�/53�#5p3C9�7�˚ſ�S2��ʽB�h�̰��4�hKfn�kR�6��x��0�%�^�!��-�V6��1��e�E�����B8/A������������J��M�:�y�M�Z����ы?�0k��ooZ�<�:� [�F�~Q5�hy��A��;�x�D�^'���P��pV��))p��`l��l��c7����0�S�錪:�8燁Zg��0Yg~�ڔ�{�L�]n�|���O��w���sηi�� &���8��F���o�m����"@��xf���sN���pcaf{�P�&L�ˮq�������''rb_�p�}.��!�9u;NXbx�憌�=��/�!�����O ;^�XUV���P��5<��SZ ���m�v�;f����Z���-�7R�'��uC&Jl@�h�T��Z� 8?��{��@�)����S�j��O�9.�<�;)Q`�@n?j��N ������w�����(xQ;���	���҂ŝ%��j��.�ZK��^���RY?M�v6%`����^�c{-ҩf9��un{]�n�� ��RW�%mJ�7X�=a���捔��E�-��τ�ƀ��������AV���Z�� �3=3[:�ưZl�AN�s�ȩp��:���X�?�Yf�`woKA*��$;p����Auh�ư�_'N8/� 2��b:�2dt�!ֲ���B��*s�O�� l{�I���j�G��y�j(M��hU�#�z~ُ)��[�����f�rR7�=ir�%|�����j���b�'�S��&��֪�r�z9�(F6Q*|�!��9���$zX3C�t�V��]U�����CK<H�N�l�K�z>��T)�s�#���ٴ��{����X�5v�	����:a�X2*7�&���E~>da�&`��tG�$y0��P���6�0BX�w�!�L��;��`�ce��1�6�;{�N!��01S��4TBS�?q3ţHq�|瞻(5do'ǌ{+�Hx"nT��R�[`��ˊ��آ�	Y�LQ.�����t?b��g�L�U�J�\� _A�b�`gل:��埽3}����}�Az{�y?S-���@<����S��nT����/���E6������A�+�p�c�}�h�/�U]k4����}�J�L�2��L{y�Dy:�JT^��h$��T(v��\�ig	�V�F,\} �i5{�.v�Y��IH�[��[Ԍ�e��OCT+�;3A���dk�W�R����'�4�5&��OM>���p�Vb
�UU����4�(��(�'�X
�_"�} ��pN3�y ����4w�����u����X4���9�4�{�{cm���#,6�(Y�HHCFw��1�ئ,��.��S�x+$�]k��_!���2�L�,	վ���ö.1�˺Vؿ�ha�E�/�c%Yz�S��^9j�6�=�V�KTP�.��qR	E�$���~�w�RI�˖_�'�B�B��/�SfBX��@|p��e�x��Uy �0�8XiI�a,Xп��?��ǁe�I/If����~����Q
�Tw�B�d��/A���/��
*/A��]Ϟ���27�r	^{Ϡķ5�k(Q9Ga���gh`UZ���o�c��-tc�����I�y��Ώ֭�*L��7UK5�T9mk��f���K�y���U7&5[�Q�EV,}��˕N��� ��@�P����fB-�(wB�hĹs�k%�e;����j��e12�F#\R�&�D����u���[�_w�0�%J%�?C���ʭ����G�Q^ih�c�J�v~��A*[8�̕�Ϋ��:�1 %`��?�ںw�^�M��Du��`&a�&��TI�с�,ow\��+����N�pEV3{8�.�z��o'k������1��85����6�_l�&�?@�|�^L��ܥ[����[2`=�Dgp�o]!��	�|�;�T2j!ј��U ��o�D��D��:J�/q��9�4E�C��d-ЂMH�ܚx�S%����w0��6$Q�zt�J�S�\=v}��~_���I?k��rh{P�,K|���%�^#��[9/U�D?�5Ot��.�Mlx�t�{��Ca�A]w�ZRW�L5{$!����	x�B.o�'�vK�����qN[�Ro�䦼>�$�WM������Zƣ��3ѷ��v�s�m�'��|�d�������qc�'��`���BY��x�a���g�wcE�Hŭ����f~*�넘)1�c�`���.�AG��/�m���H?��������'=6&�Y��H���*�\�d�.�#� �*á�eT�� 7����ˋ��@mQo�c�k�1�/Ls�i�H3����e��x�.�.H7�уݦa�V����*�~��KR�լ��J�WY�?kp/A�p{>��<��)S���u�DҞ�y�)䧋Q�pS������b����;2L�_�9�?眨��%�+�g�x�4�t��'@��G��a�C#W�������W[aj���gZ�d ��'����B%�b����i�������]*�?�7^E��qDS>O�A���
Q;U0�\R���J�ble� ����-u?��z�(�`�#��al~: (U��U@k��d�����؟�����f&Щ������e�U7��@�����t2���`��S�>>��΋B�o{"���<�v�/e���w��<�n,�q$�}�:�	��6e��W3��`i��lVOm�F��+-�olC�Y�ݷ��?��(�!)(�Z0O��D���%hjocΛ�F��ݖ�n��bJ���ti z��wP�B��F;cwp~&�LĺB��o�a�T���g���[�ڴ����هp��'�Y�Q"%T��t�M��6�3�m���*�
ū�N�I�^�sS��Xn��,�v^������N�b��m��Ȁ87Pl����	Di��7��1�-|��Hy�B��I-�VA�WA6�,��������6��J�jG@y[s���b�$�un)	X�5���
�k���`r/S�ݧ�Q�a	8, 6nb�����D�M\�^BH4-C��ا�/�ZHuW�c��f?DE��jf�C�]4�[����+"��_F�����.K5Oy�+Gp� ��M�YC}�q.�/%aأ�9�k=҈�!�w��:��E�P��a=hHnc/��i�ƙ#$$���?�@/?^�n��4���9���\9�E��.p��9�?d�jt9|��Z����:��M7Zp�)5	���nQ��gJ|���K�;� N�F������)�\h���`]"w���'oȢ��S�I��0�{qM0�{ue��*�g�E����1�"�ɢ6*fV�@rr.4˖�W�-���1Z�x��m�&}zm�K7�g��Aa�8�(y<Oֿ���]�/��7�[��m�z~#eU�d����{���O�5�l�U{�@
d�e�w�P�Nx�EJ��қF>�����
�W�i�GA;���k"'�Y��F3�A���eV}ˉ�\V�_Hw'2�"���X��I�vײv�/uH����E_B��\b>l���'�ײ�k�%$,����������ܥ�$�|ۨ�)�Z����IZ��aw�FC�S����a"ϫ��@̨�¶�x?V�k��z`�h��`YE���&Tq�p9T��DUZ1�T��s��
<��P�[�ݡzx��g�����mF������c�k]V}�=�7��K�o�@ΰ����RI[V������k}�-]�U�=z�lzZ�o��J�{U]��Dش��3H18V��np���Mǁ����b�oI�H!#�[y�B����;#�3�0"ȔXC�1������
�@0�:��肎�La
5-�8Uy�����	�0��L<��9�`�����e���Y;�;�������mk�e��O��2ȴ�y�_8�|,]��fuB)䉇��B0V�X�'�l��b�	�zP�G9���R:!G��5���#�����0�?'Q��@i���n07f.�z$3����XnƗ=���FgY�q/n���8�T�g-�Y�e�Fi�*`�����DW� �ߵ<����}
��>�N����BZ�wAU���)yc�&F\>��1�7),e�	���=#;=����:�=u�7������"`�/6��1�|�)9��,[��%җ���&�BPUmJ�X�R0�2���OVsS+����Q�LSc�?�Ȣ�!�tN�G5&��.������.��+��L���;9��5M{�m��O�I�ב^��)��hu��
���|��ؗ>��R*s�O.ߵ�8��	4�]
�Լ:C�*XvT=�C4r\ͩQ%��ń�$5a�)u�+����C���"fu�@dX�f'Iz��{/�w��Ӯ�Ķ�D�G���=C̾���vN
��U]P0�L3$k��N�O-�l� �j�_b�V�:���x831��OZ4z�t,�9m'��48AUW4������R���f����w!��J�_���ʭ'F_���:ŮF'�J����F�X����CՄPM9J�Q#,��z�A�s���ϧ�v�}�p���{Q8�!���{�t�� ��֚����^�.[5�����������#Qp}�}��&c��>��Y��fF�xݫ�.�L�nϋ/y�q�s}��֙��;m�M�S�U�E�s2w8|b�'C�h���w92;���/�؝^�όtd��.D�f����?��y���n1j�HZ�I?t1R.�
��K&M��	ט�[\��u������0�
��P��:���
�ߗ�GS�= |�q\�#1�6����k�|���F�_/�*v�D�%2Vl|7ˬ^W��(��J-u�s�?;��(
|�;�5���6q?9��l���W�L��1��+��WT����l�-\(I�i"�*w�5�̥�zj엗��ۂ��oڷk1�'c��ϹGM�:<d|.�>�ڏ%�t㔈xD��mg֡ƶ�j�c^�#}:�L*6��1pW?N,~�� S�q�B��Q���ٶCA�����X��9��d8O�\#���7�6~h�2rgߘ��W:$��,*_bi�%�v����9�v�i^]w0�b\O�i�_G���=q�q��-O�8?���bTߓ�>��IBu�SÈ9;?n��(��:]J������5>��pp�D��e�dp�@�%�	7��"�e�pm����`�#���s�����2
Q?I�!�.�D
�oh`��	� �a��~�d�h�O e�o�Ə��������p�,E\KM�T�G�f�TU�*��7椤�.W�m������L`vM*��$��/����'H�MD�v��?1�_oI=�8���E�.,�a;Ⱥq"V�����t�9&�K��	�ŧO~J��(�#�;�\�;ǅ3�D߯��7��:�Ȯ���b��u4�@|�б��퍟.��^��*�Ra(�8jM�� ׺T�g-�w���< z"�v��Q�cZ0���i�!ː ���L��Ցw$6�WT�5��y�8��.��j�|�_�dh����L	/����I%��62�� iP�	����)�o�=�G�\��J�*�ȫe
l;2����{�+�P�1�<a�q�+	�Nn�q��)(�1����V�i�5K��;�-/����Kq��| �#MyKZk��lA���'�g��0��������w��B F�kf�(ҏ���/����v�ܦ\O7�M*,q����q�M2l>�/���0���� �"q�c�����hu�X�@�,g^��POj�Sw?��h�EbL{㿙�$�4�Z�褞��-�*��OCLv���)�"��U��ǴK�9~�N�{�*���7~�xֹ�w��$���/����?��?y� �7��!xkW�*;��V���.�pt��	�0`��o{nu0���j�u��;���CJ����1�Ha%_�5���p:��CA S�:���7.� z���޹P��F��y��.�������_�5�b�ĩ|˭L�ut@w>�鑳k@��ϩA�	�( IH8���&`iY�
Ԋ��r8���h���Z&8Q�����ȩ���]u�B����l�7��ܕU���;ku����D�9Lg��7�դ�������ZX��0+~��!�<�h��Q��;�}��Vi"tJh�>����5�}e��>��WF ���a�S湓m%m���P~�]�`PN�]=��n�k7�~X�i)"|R�_ᭉ��}Z�fsy�{1�y"��,� w��w\u?J�o�}�"���@K����dF����b��v�,LbN8*�Ab�d�8���I�n�Ҝkl��W�&2�$�r�
!-,���Qh�&c-j?K�`����;BbR�D�1y���f�ǣ��5�VCdB si��|>V�K�8�:�;�I��4p�o6f�uyfd�c��m�{��\S]�tF�a:����|�"[p�=+��V|Y��yD/Op�<��ݤYM��I�T�Uu��1�������$�~�o+���IեFT��/A���u�N�I�4��T� cyM>��f��wY>���k�U�bʠ�@H1�_�ж��ۇ����\�5��t�0F闊�쓗[����`jk�������@ k0����� ����aY��;D�¶�%����-%�c��S�j$A ��M/���<�d�'���V��� ��`ve�{
��Y�/5�PJ��R�4GW="��%N�C~��T��NTs)#��l?'�$SfZ%+�N�����/s�Y�_�x3Z��6���a�3F��m�����p��?���r�͌�U`O�&"�����h���M�Qg�y��O�:G�ķ�4����z�&:��<�/}��8�e�z��MYKQ��5�
?���1�TI�>��#J��5�x�E�q�G�-Kk�H,�ŗZ^��4������dy
[W7X!%c�35��*�8�ej����*�<�ֵGy��no�l82�\ ��8�T���Ta�T�E�p�榈�i�zn���f!Yc����h��1N_*l��%�6���_�ޭ���mR?t�0a-��ES�o��C.5�|XMz�ٗA�
I�愂ra&�����[����٠��?��q���`�-����*x�5�,�/	Ă�q ��2h4��mP��14|��N�y:g?��{��\��ۀ��	#�f��+���.����=��a��3 H���+��ܖ0�O�Y����~��@�;��},
#�3|�L7(��e�~V�����0�Xɯ������bN��j��x���?u8�i$��žRp0���t	���Ƙ��
H���x)��Φ3��~`%��K�R�{�����D�^í�*!Pݼ;T&25�������j�q�
r
'N씪���7��w�ժ#�s�ʣ�[l����꾪�^�T�|IR�R�uML��������y��,n�W�&�όaʝ�XV:<6	�<KK{�V U1�4�<��'�b��TWdYu�!Wm�̃���s	�0�}����ֆ�w��70�]�4Y�Ug�A���0ۂz�a=�i�p��O�=]����O�Ճ�W;H��Ib�{�{���']��
D����FД�Xi_�Ƣ��JM�����>Eㅚ�P��j�|~��9�A3��[�/m���lӔ��i<g3}J�PE��s��.i�����k���9k$�OAHŸ\e�*L��R׹TE6�H���y�$��d��qJ�AT�r`�Ʊ8����[wi���"1�O�J�����F3ȹ4H�qm�^>|̄?cEG�,����#�#��7�Z��C݊J��(B�.d�T���K>]� �F��(*1���"dr�L`T��=������x�����'x0Bv��Ő���A=��qH�Kֵ;4�~��{S�ϳZ�"�77K4�;��ۍ�?,��&���1�k��#&	BDO1x��<�nC,?�.�Кsڍ�E.��$��yԎk���J�E�r�����YWd�7���J�����(�/�T`�6��ޜ�I}פ(�*V� ��J5��	=,Z��/��D��3�ю�{HI�#�S_E�>%%��c)����r�e�G��Ud�R}��s�(��0o�ȇZ�8"�CIK�5���Iw���2���I�� ���e.���6�,I'�8}6�!��zn�~㍍����i{m�g�:Dx�B�$�ێ���܎茓u-��C��Ws����I�S6u+��!��+(W��{'��0<	�[�Er˚$�4��� '���#T|9����p0%�w�!M�o�g�,�t	ۿ��T�|>0vM_��[n/�M"�`c3�o��Z"��{]"!�A�qީm,��4�qxiL4G��]]�Y{�NF��<���C�!��b�.5�L���{)���~xF�Gb��Oj�>��9�!����>:l��ݚH���k�/���\<$	H&������y�xF	�_�Bsc�������h���L��������������k$����iY^3�y&�;��,,)'퀗�d��D>W�`�!v�2-)X'}E��M��?�п4п��U�^��3�l���+���/x$�ꓬ���Ɏ��2%!N��a�d�g�W�n԰!H$S_��:?s-θ,H[8�0�O��4S	w�hV�2�n�1��ƾt�(4�aˈ�}�����An������t�o� W)g֠�3�Hm�-�,oc#���"�b�+S�����"H@ѯ� �ձ��B����2�nr���_����cF���$ˢEc�ʍ6�;{�)�p�QN>�Nɒ�lf�u?���E|u�\�"T�6	�0�m�%bm@�ņz}'��)]:���BJ��OJ:�8`���x��Hɪ���,y�E��Mc�U�}+����e�� ��@�t��ް	3�����X�7��j���ebS�E� (��El����������p�8B��'������d�S�!�d}�_e���:�3̉��Z��s+G�e�'7��%\~q�RB��B p}&�qF���UI�P��(���woב���+wW�A�;�Y�k=dK���Z@8�A��3��
�6�Z��{��r�6:HF瑉!���=8P%��������/ל�]�p�n�%�r�%�0rށ���2������֢�m�{;c��m\����Qp����u9B�̲O��p��ǃZh`i@�;����A���Ԅ���}��-)f)R�PpST{UAy��"~ib�Y u6(/�6���$�#���x��'�c(s�ɪ��i,��|?��R,��{��9��t��!�����G�Z�@�����.�BR0�C6]{&֥O�^��#�a��ol'���tSN��@�R
\_��P��N���j2g?�!o��.=YNq���������)[�r��Iz��%H��=��E8Aa�{xe�MPe��|᪝Xv���3F�z�@W��i�i���O���#�RZ�x�b���ߐ)/^R����:�v����;]cb���MF��*p w��g�!��W�;N� C�X+>��v��g�8e���b��N��'i��U��z��f�5��I�V_U�&��:NQ���(��F�l��/vt��[C�/�d��=g����|���`zj��W�>,=�̦ϓ� Lx��'�.?x�9�ml{'T_d ��߷�9eU���H{�}KU?x����~����<t�q���TC� [ly��1��/��h���0{��@�H�,��Tozʱ�Q���哳��FR��e��N�����Qz��a{~��j/�h��O3������,��}�2k|��/oU�W�٫!\�m\��L]���+�Vw����>�����������|�����^�o�~$D.N��;�5)��@U�6m�v�pt8��0�:���H Enƺ`g�&7뚙�&��������( ��J���~ޟ��ㅐo2�h]`��J�͂����8�>���h�ȑj��iT�@ ��Tԇ��'���V��JY��@����;_�����r���8��U���AcͰDA��ҦMM]�ۀK�oդ��ߚ�~��F�Oc�f����t<����4$��[&c��r���Y0���"]�����,]v�L��\H�buBaǂ�Ŷ��
�_�PD��czcEu��\Â�;AY�w�1S����0*��H%���5��Ψ�G�C����b=/o�7�"�P)�&��B�#XD7�E5�Ђ��up���8	�7�֕f0jx�+:xѶĹ�Ju�p5��Q���t�ty(���`B���M�:�e�-�cǭ�d����@��
&��LTAÓ���:�Aᒸ���%.ͨ����o��@4��szb�������"o��Aq�M�m)�3���)��XU�](|� �kת_�LH~�^emI�e<g������j��	�@Z�	�4�|�l�H[}��o��{��x���c�%Sº� ][KSg>7�Ɣ�^���EY���<Rr� e����2і+��������ș�ƺó������$�{�)�d���gq�Ѷ�zKr�ɝ�q������ׇ� F�:	�\�i����l�nJ�7��*&tBJ	)�:=�Id���m�BKΕ�_S�y����H�Qзl�*�
�j��V6�诗�)����.ڴ��{����v%�3�G���`��6�EC�pn�	#�UqQO��yN*���n��s|9��]�X<��Mղ��w0��p��v�$�"��'4��k$QG��e���0�v)�����I6C�M��|���́�����f�IB�%�ڛX�I]�tϲ����S��;)���N�/|���l�i�������_3i��r��M��b����@���J���i��%/ߵ����4 �� �43N��e4�
,�.�x�o�Ը�?�A�ۭ��;��)'�sW5~&lb�H>������"u�G��mKb� x��Z�j��*�ɾę��D��p5����^�fFl�%�؁�d�Mm2����g����@������+ƣ�?��.��DYW�����n9*�ҾA������'��?��Z��C�,�����\�Ju�v�����Z� ����x�M��,u-Y�UR�ؠ �6Χح�Z\?h���r��KYs�����!�=���#s����7h��&�n]��8��&മW�88�t7�b��t߱��%w���JѻAE����QQ�����?��^�D_�x�r�K.���ky'w�q��"�*���C?vS�(�]����rAP�fȚ�ԡ�܋�j�(���[r���x�\�����ߔ��o,g��0g�,�q�Tk.���zV� ۪����%_�3���c%�Ϸ���$��U�$�K �����}_QZ���R�_�AX���^�I3vVD;g�4 ]ҖO` y:�1"P�]
���Gj�5����t���Ŷ#w�<�K#ċ�9�&�N���6�<�����.�&�qG=���B8 �S`eӶ{v=`�
9��W��Y�VϰY�1(�Q@Y&�İa�J��'x�s���i��k�ĳ+Xx}���t��%DP��8QbB���l!ģH"� �����ͣ�ޝ�� ���Y¹%�'4-(���S���U�1��z"�y�@�����E�N�_d�aǸ��I΁z���M�J�K�h����J��Q��%okF�= ճ�!-�7����E:s!��<�RV~~�� F�@��gwM�杕Z�͆y5��T����h�cR�2���/V�AC�A�������ăC��J�a������ńW8A jH��%�P�7�F��ؘ]=��2��.��,7���>_�IKR2���:�u�2y;����x�:�l�)�y��W�e��O��F��΢�4�h�0�4��-�k*�O�1;a���DKs���w�d���ɚ��36Y��f��>��`���du J6{�<|65;ꑅH4P6srUm�5�*v(�/��&���:���P�� $X7�0s�@���a����G���߲�bT.ޢ������';8� �\��s�)�Ԧ���`�xK��:<��P��h���w��)��!��dt�e0��/�CfS;9�7���%	n���k���;!�am{���'��Y�HWr�#�|�ڣ����Wk��݉�o�C�l�,�qm�+��
 N���2w�k0 9C��T"x){7�-a��.*	�Z�%�*(/{�=\�b`
�$5/�.�-�s>+l>�ޅ��a�pz��]�{vڏ�4"�e�}%��C[�����J����u(7�9e�`�6���z�О�(�%ä���h{�)�+1����(�	��de�xӾ�`"^ O!���|=�k.�
ꛁ|�5��o�2���Z�zja��`s�`�M��鳾���ep�u���wu�����]L�`fd2L^���N�T�;�$"�!�S�U��������}�c��̖��1��:TML��5��@[�a����`��uDa�nT|%�[w��,6�&,l�~�|���c�JǅG?. ��ʗ"+Ud�W�<*���` *8�'�y}Aq8L��=$Hv�\D�<1�����;	�e4_�e=�|�������f�[�ur�*�D5a�%�J"�,��\)>�R�(����[�j�6���iط#G�<;�D��L�X�T����q����yl��L�z�l��Ҍ�ϡ �bD���l�h�������!+,h��~��q��F8�?��9���/�5�Rs�1���E���K"4���W�zA"����Tu�ఋVuPW%�ߎD���{t�� pߡ��f��=��F�qѠ�^�����<�Dߍ(E��0qӘ$�j4��e�n�D_4��P�ZS���G��-E��Ź\&�����*��O��߅Sbd�S?�J�r��l���#�/M.:��)�N*��3a�W`j�]i�ɺ���ǝ����yHTe	��[
�Fy�b�:���?'\�
�8��u�]�cx�&�*=��Y"���<F�Ģ���ݤ���v��{��/b�.�!�o�2̆�K���=����f���^�u۬КK� �ZO�P�8�:j��� f������PW�Ӓ�09!94VĊs߮R">�� l���r�f� ����/i��wQf
��9������m��%���h5�$O���C�P~�3��.w#r�;���^��'\�} ��kN�Sϒ!0x��,�o��S�~�e1��� pw�58u��:������
�
\�7�����D�;�V����#�dվ��9��`�Fw��dΤϯ�x�(�����T�����7C
|�/��|���w�7�-����E��
�Id^�l��}�{U#r�/���´��=������ݙ�HQfl��CQ�Q����8�h�SZ�AHC�b����2</�1Ps��x.`4�i���ţ߶�������%L�,���6t��T�Tt����K�t�9ui�dgg&:��:{�*��5���4�޳"G:[.��Ϻ�d����%��7@�e�_'Fvi�#T��D&�3�Ѣ�θ�R
I�	] �3R=FZ�U�9�14N�|.~���YǕ�Q�>���aRt> @��P5'Iڃ�����N���ه{1A|��w<��R��X��UY�q�tl�[5�;�y57��D+���P�C�n9aFS0B�l����@-�y�I*��Y������r�*�2��4�X�%ԃ^��:z��1�ޤ2<�!n��Oy�������0��A��'Q�����¾��"�,����o�w26�(Փ甙�Q��f�����y��
��Ʊ��@�P�6�����e6����~������ET�,���r�ʕ�[d{�uuo"�	O���+c(8�"�rmO2T���Cv*#�w��:�&!���_p$����{t� �� ���8�!^�rz�D�R�*�(0s;b������i-�#���L��4�83�uI�Ź��``͔�3�_��V�_K�SGj̧���<�f�4��I>\ҐŜ������vt*�N�F�`�qG���-���=Emv�	����7L��R�&��p:^?�M0���%���$CC��=�-!���튳A�M��
a��9���(Y,�?F6�d8;i�Lm�j}�`����U��X�_�l;ܞ�e#B�q`�׭s����D��"��JE��k��5)��D�\�3��o��&%o���/�� r ��n���� Z��U��.\����#�`������,�#���q��9��8g���ȶNubA	Z��O��{-hY_?`�h�8>o)�N��[�U�6�n����==�#�W��n�p3��r62�����?;�N�l�煷`��:%E��� ][Ӝ�Ǿ(��O��L"�P���pͫ��]V�D�����a�Q$q��[�E�c������X1�ͺ~���v)?�`49�c��Q�W�\���|5���Cd�P�%P�P�A�{�Q�d+5@���v�Ήo���z�=��BF�<��)q�B�i$6 Ь��;`L�jKxAN9�gtQ��O;�����\�TfIy�N�Nw���lWxj���j1�^p��������E�ߑr?���}")�Z���n��#Gsp����R�=^��8�ug�s���0�/N�D$��!w�=�قdȯ�F%�B&��>�u�_�l�F_=���O�'���f�e�rE6�>+������	���@�I侀(��Y|ӣI2�g���ގ�rOؗӅ����G�%-��|f�\�,��@�� 乗3�c� &�)"��J�H���MW���r�j2��e��/1�N�Uؖ��<J�({��I�P��L��d8�|�0���ħ�zz�9�X����>��[=KcM�m�g�v�b����?�l'wZ�������۽�E������&���LOh0"���;ai|Ԧ��ˎ����H&�n�ı��vU>v=W�� N-�����
�|?:���xw�X����}��a,]�T�۸�K<����v��H�@�ҁ��= �̑T�m9i��#�Α�1BP��6<�}S��^����p��iǎ]�܏`t5�[�GU���+/TB1=�&����#� ��9�`}]��G�#b���+}
�l�aCB�&^;����Ke�,@�}'����de�︔���'f=��0O�j��JgC8�]<�������~�)3_���=L� H�/��B��X4�L\.�W�d~�����Ü�RT�
�0��v�Mi`��B������-]��bH�#��#!�Ȳ�f�64�ԳMt��&&qp�e��Hr�k�I��=�m�cQ�Ѐ o�P�<tc�S�p��	�	65�g>u�]�G�v��XK���r�v�)�	~��S���fkX�%��{+���HQZ�=�֛YK�^�܀3LS\oF�[}+y|��y��6���X�`���|���p���t�7PkP욄��_��~u�vFUjG��6�4�@�$�-hC-�^yX��5e׫��yC{�{?�����t����Ro¼��
�D��)�vgd
��"]ӀbW%R��7�`�\�S��\[��hC��V_<_�
Ia�9��`����C���7�"\C�n�Ќ����RVo���I)XI�� z�N5�8J��P�ń:�B'v��:�,�a��+	�k�
��dm�d��uF+���^5p�Z�����7h����~��c�Hq�XR�paC�<@���O��B�	SWߔK�y����k�]+���-=�ع4�s��B�X�7]��g�[Z����X"���WH4�V�ԧ���_ 18:�)mz BNI!�����x��$R�K�}�L� �p�pح��|���ܚ�'
1[�)���&~`,�9�_�s�<Pjv1��S�dC\2Lg������-�61:��>S�t�4���m�/p��E��{O��d��3�E���E�r���G���s����w��=+?���#66�X�~���q���e.']���m��t��:�Sot4��/^@��"��S�2�egLz#��6��J=o�uu��-\�tG�>EP�̡�{c��6��
E;4�ŹYgfAeA1d�CXIS3��o�Κ�X?h����}o?e�$B��Y��v��É4�eVNax}�ư��c�N��S�SH��ΡsE�[2��ӓ�su]�(dh�<	�`�����q��"�u�l�@��)�V�N^�$=zg?/�/U���M&�$�"��e�Zlk`�r�e�є���ɚI-r�.(��N��ѳ���j�;��<)6��SjK�ů��y���_����� Ȗ�y#e��=�-I��Y��cN���s�{��Q]{��*�\�.�&��4{^�W��*�����5K���e��g1���)������['����Ҕ\Z!�ք#���4�v;������!�� L��0���_$���f���ڪJ06��`�,���_pb�h>4cU�z�j����`�m�R"�6ob �r\��rI���*� ��ȾH��y?[H�_i� �n��|V��j�j��EH�A���Iȫ�)���K�=
���\+Uc�vHǮ��>�*��7^K{K��4;1s���x����҃s�ji'�/�.��/��e٭���s��;�ҘA�LA�V&�7�ӓ�w��� 2���Ү��Y��e�#""ܩm �e�c�K� u蕕�`��v����zKc���� 	n����.�u�)nIX��N��3�~w��9F��⎕7����xn�(�{&|���_������\���h��Ӱ{d:1�_� M3ec.�#'��r��朌�L/]p�h��U>�RxɊ�5F���?��țؽ��8"ܳ�+����Z���Ǡ,����3�	���5� �ŗg����J�N��M�`��?]8S�G~�|�.�x_��=��9F�:[��}^�H+�[��|oSܲwg_@�!��d�1���
����-jn�UZ+��{���m�%�:Ѐ���8�v+�eu�ۙ���mL�����=�1��B�%'r������A�q~ry���cr�[s@M����Cnr�f��H<���4���=�^�|���Z�{[��Ԧ+G���}p���u�Lj%bC8��V\�����8���h�f��Z�Fvʽ�d<�xz��j� \V����o셀�S��S��o ���o���S�А$Y��0J�̽�������db������x��(���T������ӯ$ `9�UM����(%�.F���̳�&\JQ�Պ��nu_�פ���a�MJf�9�9�r4��	)����8XK�j�Y�� ���;t��p2�+��E��zb,�S���r�u��/� �CAq5u�P
-��KN��P��fX��#���9[�� ȱ�*ϓKDx�L�c�z�RX�L���� ��r��쬨���G�]�Y
�^Xc�]� 榻�eJqI'I�>o��O:�0��f �4'�&�>8�e�%; �?���H���n���ˮ^��t��j�]��=��aӔ�� �ߩ�7�ݠ���!J\9�A))1����O�VX�;�gC1We��B㕧(/-$�uxQ45 P�Yq�H���d�J�h�N`���,��&��'r�+�0�P�
Q-����#��J?����P�W��@h;��O*�>]�c����"�����a�	�~�S]��z�[s�V4I�F��&�5 8�X�B�!�줥��pL�Y*z��!	1�~=�@#h����m՝�*d�؏��^g-/���FR��~��+#���u��~%~�`��C���W�� &���}�����������5B�sG�䡵Dg��Y�nX/獣t/���c�j��q+�.�+ [8x� ��z��z��r+Eo�fw���D�(�E���s��]�qj�kNƮ�;Ճ�������ՔH�#���*,z&l"�H���Zi���}A�ܩ�N?9��ؠ��$Bچ�aR�VL�L�aN�b����Fr+IP�i�L�ܵ	�(��s����&Q�Q��Nm�l;�z�B�J�̻�/z��\�v��7 2R�	�{�<:r4���͎�è���_������|�6X���5��F&,���2_�6`խg�q���
�-$fzT��9Мy���1�?Eb�*L�ٓm?b�J8�tDi�[#�4Ǌ�g������x�ʉ$l.m����9b$��B��t�h�R��N��8�	ρ�6��N}�Z,K���h}ws|��qک�w�S5I_`!s utX'�1����T0��q�"w3�+D�K�8:�:�Ǖ�І�_��l�?xqj�V�6�}S8�Ƿ��:�.��Vj0N/x�ZM8KjG8<\��a땨���[�j<K�|{Z�������<9��Ŵ%�rSM���+���S�w�lƐY�2mw�s��]��:�n*���N��l�ein)W�è G�Ai���q��oT{W~��o%���,���wx�X0x�n��v�4�j����b�)o_m������;BA���G1��W|Q���&B,�l,�3K��B��)-3��)f����g��A�;�f,����w ��3kV_pP9o��v{��#�ũ����x�?��'t4#fF&\�g�E�._�f�KH���}�A�l�:a��yB�
��h�	R�ϖ\F�}OnW�Ҷ7�
s�U����A��
�e�V"�rS_ʨ���9��J��\9��)�O8��'E�z�S�J��/�f�k��A����ͫq��y0}�2�X~/]7^��@�}����{u�]���.6ȓN�6| @��&'K�Z�οF2$���}2��!d{5��xA�o�"��b�:�6�C^�l{�¸,�c`�>RtZ�\]�ؼ��tM��H��<S��V�
�� ^���]-�'���Vcӭ��chQ�grjc{��k	o�˃M�
S�s][�Cy�nqX��}oaN����qR�!/�n�Ǒ��/��+������I��}m��Ʀ�M��/�2t⼪�l��c�8�I�3N{�l���� VF��Y^��M�Kk���-���1�oQ�F� ��.�>�&����E^_\ �T�H�@Ԇ���˦�C���@�Ǥ��J��G��ƭ4��
k��ǔ"$��Y�d��~�lnh�rw���Ψ&_�<#O�FAU@΃^+;EF���"Q����03�:�t������J}���YK�c&3zqۛܰ�)c�x�JQ2
��OH��`�1I���k?��p�cx�`���i�{�'��9����Z�ӵ�(
o���tN+ÜX�7t�	2�F��-�+��^�Q�=�Z�EI��1pn�h�ڮ�e��p�Z�6�5��*��@h"�jvQ���*Ҁ��?���3��r�C� ��a�Y8�̓T^p�B����a����;�/�7cAO�YLH�~�U�/lM�Π�(��~.)
`Jn�w���hOw# �ܙh!��f9���x�o�p9��"1�����=	�D(b��&��)�r\��t�'u�'�������&��:C<�}}�%�IXٟւ+�1B�=:�)��:M��呂O�@2�&>B�8�R��eι�6��7%#�x�7ΰ:����#z�z��6��6�1g{]����	�ܫ�|*�w���|T��h$
�.7mz��!P+�̪;���|qޱ��Ȱ�SR7���f�W0��p5��1�_��{��ϩ7�]���7_�[��˰$q��=S���59 �?N(nՔM[h�/x�[��/��M�a��jK[N��Kƛ�'L�[�M��wPJ^�Hv�V��-=i����E�����T����ƭ|KātW���
�����r�J�6J���2�Tl~��)=I[�6B���D���ٵ��q�S��y<��ku��4��(
I��t��Sg�".-����+$�z����6�LD���S���F�@u |�(o8��NB�C��
v���T�]�Y�Q�\٣1�TOl)�[a�3��)�|_�/X�q��F�p|�?2Vx[��Mf���3�x�k̂��1�c�7�V��®�}P�A1
�?����L���4s�r���e����8i���� VV����H]��N��n7��:_t�
� 60���&�;Y>S;<����Y��C;��Z(�Ý�to._ԦC��n�C��h���mU#Z �V^����"�_gk�꒿����e�c�,.I$�*%�����j4�R^~9�h���K��ΕΝ�<ey�����6�p��oҩ�L,�[�h2���G��zz�!�L�a�v����i�ː��6�1"�|?d�Ʋ��|����3�����_)����NCuY��zϏ���-��o��&á�B��~�h�ϼ"��Ј��Ԟ &�
w������yM0����Ak �v��$��:�\��vq�R&�&��kM���n*0/�K^���N�x`��8`��/����%ݩZ'�D$i��ܾ���Ȯ��\�樂�F�M�%����#��R��	0��2d���+�aU@M��3�9����o} ��7��: ��L�ѩ	�'Z�.QbY������!\������/ib2���� 
v���d�=m��Rɲ��Z�v���;ްT�l��Ԥ��Nӗ&]r�b�[,�u�=Ȝ:N��k�Ri�寮�3a�p�;��➳=��Eb�-�C.�1�0�_%�UjA��i�j�1��5ƵS�D���<z����!��A΍nz�o"�2K��#06A������ܶ�R@Ba�o��d�@������ei˥/qcly�O�FUz�ܑ7��T5pa���ڿ�U�'	�|�RT�<q�t�$M�S��Ѧ�`��є4 x_��fMu|Oӵ�K"=�K�f2F���K3�95P�n$N_&,A�ЧL��
w8�?��9Ξ3�)��1ĭ��Q����jA� ���[ �e{��e8Nr���M��:C�@v�la =u``H.G�.Os��.B{��Ё����b+��ׇC��-7�k�����<�ظ:,tw�n��OL����ނ_� ��1�(�gΓ�ї3~)w��1]��rT�x��p��Q�u��h���xa@��O�ۈ�tρmao?�3�,�h5�7D�&W9T����g1���N�.���+|!��d$���0<���Ů�`������X��%��3_h��R,�O�_��Yܣ�E�L��L ��ӑ6���P�A�D��xж`qC�!���/��/��s�5M
^:7t�b���gF���%��'VX��c�[ݫ3l[
 N=���n�PQޕi�_��Ф����eΥ{�Jd�I�F�[���L��us9Nlv7Jc�Q�F���}�ۻ�zS���7�d�.�^🁵܇S\J��� |ۘ�hМX��Vl@�C���h�m��}��%���=�φ�O�5�`Lr��BR�s28���j�0KT�,��E�kxh��%�;3�a�?՚��D�ڵ��&����ll������g�ʸ�������*�b(]�5�����\���B�k�G�;�����b)�=V�L�����zHx]����5ONPN�ք��������U��1�(Yb�vX/�
A-�KD�/p����pﱹ�z��l��ÕOk��4v�8�@Y��	�ɋ}���^���"
���t������:8`��$ґ�ү���&y�Ƕ
����Sr��&���Tr-��3�w��T`ܴ��gp�d�u���������+<�U@�}&d�̰8[��}<Ê��"�������o׮�L����"k�p��?b���A�p�����ڲ��	�M�Ͷ<({�[B��Xg�T'[�45�5:�M>��M�F�Q�Ι��ӑ,ĉ���p��s�I�1�����gi�%�H�y�fK7����Ż�Rp�~-�ٺe�(��̂���2���O�4���������ܡ���:�Q7��p�X�	+'.x�%��uҚ���7�{^{��v���~f�GTb֔�ur|慄��_�{C
�QV��H��q���p��!+1��Կ೧ ��:�$<G�NC&�%���k��h盌�����p�
:N9�����!C����n�����a�q휜�K}�/H��y�x��lI����!T
�T=x���N�*q�@0t�])T�[��,(o�����e��Ty�XP�~�Lz��X���}e�gC�A`\�S�\Y����Z���%��7%�TRa+�֑�B-kA���-���boYy-���c����z"e#���\�Zf&�4�,���� ��U���`���s���F�-���e=��~n��bnD�O\R�үw?I9��e��m��d�Ihُܐ�-U�o��o�޴hE���ߧ�9ۥux�(�5��ٽ�˷�vm�Q� S��*�xo��-i��+}2��Iĝ�VCZ^X��j^���v���~׍4q#���N�̗���::�
6�D���H�p�:�Fo��_�s�@���������ALt�%�!��Y�����֟�t�R�Gf�ߝo%����Ϩ�5����M���z��ۥ�ῆ�rH�	t����g&vϕbX-VS����v(h�q����Ti�6-�+G��2��R�#����0[�db=FpЩ��T�M�������cP�u����p�I��1EԾ����ǀ[ݶ}�!�B�m��tc��b{�Ӌ21�D����i#���Rf�	��Ʋ/>��Z�iw���IuLY��Q��z�i�\i�=.�<^���i�5|�`��Q^\%�҉;7mʾ�,�	���ì�p�|��� ʢ>���&ZS�l��=�J�(Z��U&bQ��!���7��-yRu��f�ӿrO���\��N�O<�B�Pj�;����Sr��׼��`k7�	f�2fK�g]3h����Z��S��`f�u��%B0��JmEh�_��H�&���օ-���(����!�/��8^��,�����!����f��4�atA\N8w:�=��zII@w �Q5��xX�Л�ϩ8S>���c+0���@$�'�����(��E3�r�`�Kh��v�i��t}��,��L���
Fn'�{]7i@�@��m����T��g�Vs��]��U�����<ZWw�6��˞0�O⽉Ax�R���,�z*�na�s��t�a������An���khhGu���ꐗVإ�T�����Փa��団PL�:����h�(�F���eg��z�c����%u� 8�1�v:���������8�
���5�[:�	s�ʸE�E���!Vq�@Y�E��|�6�E�Z���������n�y��D�˭OI	��w+��o���o`,^��jx�;mR_d��Î�)#�7L�U�轿<�-��@��v������\�r����;�76F�C#R8$_Rt�dh�O�Ǘ�ɢ��(,�]_ﻟn�mt�x�Tx�q[g��^j0lGlv-�	NʈCt���g�t4���,	����=eg�0&dT�t"�J�� �_�Ͱ�'�qH�9D�M1���|R���4!4p����yQ�L2�[|��[�se���}.�n����1�6�7�1�4��>O���%��E��ȅ��|{
 �
��%j]X�E)9Q^�6� &�W�\-2z}=��C�h����
d�PNv��5}�0�#豫�:Q�5�5�C(�|R�[���9��Cf�|V�+gϛ�J�Axc���0V5�V�������ku�ޅ�͊�o���1�,|A����E펴���nz�͝��2��}WU�R%/X�?͟n��%�7ܓ+}wS���k���BJ�b�8L���F�Vډf�}�vN�^ri�ܻ�T��ۮ�cEP��8�����ZY���wqx*}Xay\	��Un���=����f7>�8�@��tЮ�� }�R�#�Su�T�P˒u���"����n��$%�����aX�M�`��dȊH%'H�0�?���3b*Rc�����^L�Ϡ3N��~+��q���	c<�OmP���i�o�HT�gcm����xY%���Hh�$.��g$� �K���Α�cyi�}�����j��e��Se=��b�yb����Î&	J�v�֋�t�V#�lB����F]Q�Lzm�irЌ�%�њ�c�)g+N�D�������.��Y7��L�`L���~!@� $Ki��5��n�mS?$q*!�B/B��࡭�1.	dZ�qԗ��BtUV���]����3:�T��h&4��HX��:[j�snfDťݬ��,���Y�/�J/���v���L����&�p"��]Ń�~���Wf%aY�QeE;f�Ӹ��<6U�ֽ�zz���)�r-�]�Tb�#ˢ)��#����ecz�Q�齜��3��J��I�(}�����O2���<�Fŉ�	>�ҷ�FT_/���M��
�)_
�-��m\~5'΃6�G�j*t��HRްc��@�u_q�.Zn��'+SS��f�)�����01M�G�x���]�r�Rn��LD���I��x��B�M���d��u%�;A�i�>�������enP�y����j`жv&�?1���kjX�8��S�i�hl�XJ�c�
�={�6^�U�ݷC�q=�qz���q\4�ˣ>B��&��krL	,�G�����z��{L)��\���f�lʞ����F�E�u$ВD��l�lq����m��r�Ǿ<r���:|>�gC��r��WҸ"�9a����V6J$J��?|�OL�ծ�Pm_O
(�,�p�*������ʡ8\9��Q�L�͜���\:�(P���.�h���ig��w#��
F�����1A�ajQ4ؐ�Х��2�\��
Z֛�ՁTy|���C�k�>3F��h��Z��"�qƥ/s%YN� �]y!�ώ���m�ׁ/�d�u�ڴ"�3�)O�{�ȿB�'gA�@��� ��'�-��-�Cbx������$2_�T���~��a�W\	 �
Jm*����q�fi5Z�f�ކ��Uo8I�)�_�,�Ɍ�b�TPO��-6�Z4(�`��tԉ�	S��y��\.���Fv,24�>ն�2�9c�qA\% �Cp���<�/?n�?�Ǹۛ$��p��推�T��s�k���(b�Of9��&&�1��eNT�<�'[pq�Z?��/�9F0�n��bp�3���+��-Xӛ��SyȨb�S9��9�؞�K!T؎~�
Vl���9jW���+U$���`4��1�Ӧ��ڷe��R `\s���Q,E����i|=7�6Y&��S˾l��!���7��"**�xo걌S�%vd�,�6�`�Y��S�D��#G�n�78�k��*��x�[4�ά�2�G9�O�Ff/6G1H��ۘY���0��qzPmf�`�y�:��z�Y�(����W�F!ĸ�6�?���ُ̍wN}S[ص|Y��7�C�1�~#8�0��Q\Bz�Dќ�ޞ� ���w5@�/�
Pi-y�&��ϼ�{\����<+A��	]�xq���ٱ0��&\��6�UV��t[K��N*ğYx��PT�&F�����}h<[�G>r���G<B���|yt�N�߮`���U��	C�9}�)�t�k����hX����/C��r2��j^-��cœ#�zh�.�g2+�_���Z�Hmv,�ΐ�Pg6J��g\��|+��A�@9�������|�	�F�R{t���x	#	�+���q��T���/8�S3�J �]"<¼/K"��6�`�w6h���~�d���gvլ_�l^7QL\��B+נ��2E?n�k*�V�������!��t*����B��6<���(�F�������/��k�SDZ�3Ku.�Sԡ�=V6=y 8w���9j^v2�����5l�ʰ����?�\�2SW�{��Ȋ�Y4W�K��df���}Ujʅ�=������s����	y�U�@JφC�N6m��&?���͑ú�����ZQ.z���R��̀�hB�֗ΊR�ǈu�ܽ~�#�̷"�VA/�����C���^\�i�M&�QY�͍9�gs(+ݏ=��F3�!zڊ��'��Ԍ����_H�c���+/�}ά�DK�W`ȟ̗�bX��/NO0�����Nv*S�z] ij��8��Tf-1�����1�*�� ��b��)Z�d!��E���4�)�|Bb��ɪ��p�r[�������i��ѭm��Gc!1���}���<�Ծ��ŕ%��2M�r��}&l؎��T�u���b^k/r"�\�g0HjM:d�E��%Qp*x��n�͂[��t?���|o��yE��٘W&v��N�=��:���������A��q�j?�wfdٙO��1��T�ROh��.�ibld*:�W��]��M"n�bQ}ڡ&%�=fq|��>�c1H��P�4���M�z�SI�d��/W�P����bJVΒ��QU��D�=�)1�s�l/��W���6`vX��f���]"�H���+��+�@BV�U�\=�S����\�)�0�
MX�D�7g�O,!e��;��� �锩HV9�C@��(�<��Kf(=��ܼ_l`܌�"���q�E�=�y�u`C����b߶����$�xm���V�r�M��i�_ɒ��	CS����V3+�_Q�j�:#�D��kz�����S���L� �;[W�l��ZQ�L0�~��A_��-����"��:�D����EA"���f<�'O�YmSK�\r�b,΀h3��HD��
УJ�g��EPo"/�7\Ef���TS-��⼎� �Cٚ�M �@��A�aK/B���-hk�� ��D/^lj��xw#�{fhctG߸(B�hL��$S����$��V%��%���|k��i����E�
~�!�:����S↴�/�yX�q4�49M�ݓ6���X�f`��0Z���(t�&�׫���L2u�](�G��c���$[�d�/����p{;-˫R��Hw��T9
���M����i�AeRO�A2Ä1 �T�mp�ETO�Γ�Y�]�0��/�l'��-$V ^c
��, ���W�!W&����!`�Bn������P�����k��v=�'Dce��,:��L�K8�N۫S��i���MQ=yd���g1�n^�$���֯[��ũ�p3� ��)�*��s�='8y�p	�Zܘ�e� \�P,�#�p�����/���{��S�i�\�⼎&�b�"ۊ&�9�(Y�ȅ�^�m1 g�Bq7ힰ�FAQ�Z�@�U�Mp�+@�U�{�Ҭ8;3	��W[�ȯfi*�'��s�4��4>?�^��=���e�.)qh�t���=��f&QE�_�#eh";(z��+.]Q��5��p<�.�6�07����~��%�PO�.>2d�}�+����P�>�됝Y���*��`&�ϝ��t����wih�y�my�=W �gu�3�s�3�\�غ�h�����=�Ej���e1�d��� D6��M1A0:2U��&.��o��[̑� �(�Z�Ï�L�S�T>��M��B���U*�@=1�Ψ�|�jH����L~j5B˅;��1HCc�@��_�!/��	@��C�d$�1�I���ĕeP�k[u�L���c|�'�ɏ�+"��R�D��G
D�B�Q=��� [>��Q�k�8�����"�ch1�(��}��X��bQy� ��hϥ�)��%ױ$5K:��BR8����c,=�=N��7<m\���v�W�ђN��r��S�`�c�%]D�ڂ8�U���Z�$�j�����E��������_��9�q����*���I3��TdK�y�1w�����p	1�����Ge���s^l���|02�hj�D�Yd�P>����}�Ӳ���!�ĪժQ�чm	J�F�Q�����e��ϭ�}��Vk����!F��e��g��]�
; �����<�h#J
��Ef�HC`���'�8z����6�g��׵/T?VhJ�� �n����	,�u��S�S�xRL�)��K�����iI���L���͈f���)�O�AO��J�m�b`uV���<�`��ٖ�MR�����MP�M�����j#��ѕ��
�	�0$��+�t�S��lڲ+�A9	����W�]��
F���SV�22�0?�E��$u%�'5sl{V+*��cZ{|~�dX�7�tP�˴�Mlځ��j�f�I��C� /����V�X��~3Ŏ%��E_�E�1�Z>}Ey�F� \�6�%[��k��<o��4A����d���B�ݝo�=Ը��n���,$L�R�}ދt��˟+`�k��y���8m��!Bm���##%0�A�;Zͱ���I�]���s>~-d#ϣ�-?�*�5�6���4��X��*�����"�$��d��^����}�A����E�&�(&b�C7GJsO �tR[�����0jL���>I!K4ؗ~���o]��Aq�>�XH��lw�;<M�Վ��<:����U�!���0�V�c�:x��ѩ���ihhv0�Iw���W���f�Fq`�
��Z6����1�����\���}g7r�Q)���z�z��Z�i�U]C���Y�b���~��G��� �c�+����� ��P�!~���u�3b�C��k.�T�Eu�Q�'ی��ㅹf��W�冞?oBv��n�f��l�a�'-���p&�@vl&�A"�1Fg3��QP��x�2���?C�	���ɋd�a���I`��ȯ����f%H��a/W�I����	B�$�׃l@dA'�p�.=B7<��<T���n��dF;�Do#b���I��(݁k�h`���+�`�j�O�>�MV6�l����Qb��t&A{�w���}�Á;��/�*�@-�XI=@C��@@/�$��S���d�4T��$�3�A�\}�{`B㓴ج)6����/�X:�K=Wa	��?8�ɮ�-Ւ���=��v>4�B�h,/��	 Ě�+}�i�V�.���Un4$8��~�T�y�wg�2=��{Na4I��|�3R_�+��;%(�6O�[$s�^m����?FG?�M� ?ށ���ͭ����eU,4�/���l4Y�jܹp�	��ؾ�BX&�l���r�*k���<�m���v ��"����F@��hVs�L��Q��%� ����~�_����/;]D���po�Ҵ7F���fW�8��\��a"����FIƫ������Q�]�y�K�A���;.�v��\8 ��d�a�4.�	H{����r?�X��|Z.��q�/&~�E�tƬ!��b��B'��P�o<3�����I��Ҽ��1 �u����p�~�!ǎ�s.���7�p���޵�����*�.�5P�j:c�yg���+\M�/�K�h����$zb����R��������˰TԎ��X�b]TuQ���Z%��vp�a��P܏�7,λ�����1tn*Ğ�|h/��I>++ao'��軚�S@���B��n���;�Nqڊ�/�<]
��A'#�J���d���Th�Ǚ(���s�H�W���>��C�a.��A�y!������OP�L���<��!ؘ�
t=�Hڷ��0��Z�x]�
;�Do1�<�s ^�?��Zu�5Y� 8-:���c�*��K&��X�Qm��;�5G]%���^.Ƞ	J���+D5���H�=��2MJ.�W��,�G��b�[Hz��Tb-#W'axhM/�Uj���]p��Qf`<�s`OQ>�5���z��W�� x���@�o��؟{��L��������MM�UQ(T�$~��{������iA�4Tt����P��WM{�e�Q�^�
g��Ȧ1���;d��>�A]�ݡq�ujv�uf� -&�K�)�B����G�_�׋�Z�N��'��Q�"��Lex��5�Lŀ~H4�i� �}gx��"K[c𗉄�<�u��Q�!\W螸[����i��p�!�]��b4�� �3����_����z"�z����`�X���_x�U�
}Xƕ��4�6w����o�)��4FA�?���7���~�SD�5�U�S;�t@L�!��/]괥,�P^��?Sў9�;��P=�yǅ�8{��E�t U�;�[�ÄB�~���.2t������_��V�A��#��w���03'�^�di���Q&֋�p�bݳ:�ʐ�\
'��A>�ފ_b�<�I����u���b��LO����]���hc\�2oW��(���h*k�H�z���T/��@�Zg�F0i��5�q_�N��o�Il��H';t������I�I|�P��`�m�!���y���o���I{�ttQ�!|R.�M|�I1��oKB��y`��|%	����e68�'7��Tr1ł�Ee�a��Y������fϯ�/Q6�;�Ƅ?ޚ��2��K����	i�LT��]�o���&-X�6���m"��%�Di{�[��d�.	�c%Qע����h�x*��6
��&��Վ3`��u�����
��5/�����'lQer�H�o�����[�%�C�vY�[��y� ��:��r��/qg7[�>���7��Պè���)ԩ6$d�c󻣴�r�8z����F�ܴ�b��_� ����I���F��H�=�Ӌ�G?�iv�Վ��s�Y�A�OX4c���A@,���pWF/y>��P<^Ƙ��\1a�����-y�*����"17��c��0�?ؒх�_�gI��6�P�9U�W���xbn������Y��7�ٻ�3�"��r%g�o&t��m���c?'ʷ�R���JV��)�:/���s��]�D��i��_/�Tp��S���B(�FgV��CdS���<��ܘ{�౴Đ��jTd�ł�l�%�����@8�Q�۳^k�	AD1����n/��빼-ҙ(��l���`dy���]>F����<�C}"�ӊ�����zs�d��WR��W�9�d��k�"��j�ի�#�\�Vh|_���»���[�uv�x��?�d*S�j�T�,j(���&>_�ũ�=^�{�5�nz��p#@�%KV{X���

��I�%˸�#��j�����C��p�@<��c.�k���#2<�?�W ������;�-���څ���\�/���aw��|����/-���0!.�>��k؟�0c5 ��2ul�n�=t�S���V��_��'i/�.	nH<w���q�V́?���ߚ��{$�H�b?D"b��X,kjDu�P�_)���%g����ވ
E��`#��.=
U�x�g�����VDNh��˚^�{iz4���k�<6
i��R�*aa�P��nX��|{�!ʵ�D�?�~ߗ�ی�s��SvCC҈��ҷb�����(=@��:+D�t-�)�u��2�t�#&��rY`��Rٹ�
���"�݋�����k����*j�$�-��l�����ĳ�GY<](���$��N��M�Z����9�Wz�!k3��-S#�il,�̽���Dra��V�N�-��
̙`��J§APV�f,��J�
���"��;|q���(�9����~�^��Z�[2"|�q�z�.��L;�ޮs�JP����'<IïD��l��׽�1���i<�a�s�����F�8$�5nؑɄȅMSe�c��٢a{z�?�䴠��>��P�:����G!�_�V��;B��Lljӈcjm�ĥJg��8KGn�K,B���-��[nH��ˎz=�
V��]���C�4���iҥw���:$Q_�2"������*����Hl�H}�����'|pP?�W�?��o���ŋ2JA�j��m��R;�������Y�k���j�%�o�mUt�
b���G7�jE/=����ߎ���ςÝ�#�)Q}�2a� [Ò�Rv1lI�����ӿEHR.>p~$����U��*�V���R�q��_<3|�~��0W�z�
��ᐸ�E�jLxj����@����yW���(=BZ��Ne�o\&����8����==�?uw8�iC�C���<�i]B��ig�xkM��r�.EZK�qM������{��j�#�7�e_ѳ�仢��k<"6�%�k��Z19b�}��7ƼD�Mo����gCY�X��\A��^]\@�7M���Ƞ�g��`���c���[X�VĎ�6�tB8�_:I�@k��=;���	e�F(�"�d1�����Q	�rx��e�Rn�A���<Bw��`�M1�W�ը�'�}\�6�܏�v*�w�����NA ��h>_g!�e��{Y ď8*;��.�ZFI�%��
^sk*d��A�i�D����et���6��S�U�����m�i���$��t=�dT����NOG�C��H;i9䟁��H�{�j�nr�lu��<H[+a�S��KcmX�eH0�z��!��C�F�c���iQ�`z���ſ��q ���tfZ6���Fh����3L�<n�Ʉ�%x�9�����ts,`���TʦF�_���X�3��������_#W&�\�\�׊B�����.�N3&bE��X���d��u�,���>��H�!mE����
���r�u�aЮ�;��q1�KL�gg�-�s�K�;H���qb{7�)/�P���M�+�K��.�Q�C]�W�nR�/(!��f�����?0~n�:��9WN����s�6���P����Gi�OY/dЎ�����U�h��z�إ�G]�L��O��D`$�o�D�nr���;������x���2[��sklӏ�����w��6�be|_�m���_��s'hY�=�I?&F�敍B0�2l�YKU�!+���h<cSk
���c�k�֋G���������J�s���14@����
�����$5�^e}O��q����~����Je`���!����x���~3���s�|�_a��P^��������L��o�`��D�/�$�$�a��j�~����U��D~��)��F�5�H���O=n�{�痢U�6KN����j��`8�]�¼�T܄$�#'��=�U�'C��M��kޭ���� �m����K3��#��C�I ����n��rF��E�_�ڟ>�=e%�|���w����AMg>-l�iC�V?1���	�� ��,$J*��EV��^yA����V�U��<*U�n��	y�C��.E��F�Q&�ն�n+���U�wh��� ���>e�m]ţ�F6#^��B?������A�$![�[�s�u�~���X�������5�]=O�1FgҾ����%'�#�Ɏ*|�1��!g�4��/����s�s4���h'���7/5ڵw 0=;3[��c4�������Z\+�
��0�O|.�Z�/��x��NM0}}
-:i��Ot/` �ҴS��*	�W��������E���'�f��j��\�{Ż�fZ,ˆ-�l�s
���{�ݚ$��ceն�S��.a@7�$u�ZE�<�,�z3ψ�kh":1��mAž��V�$�8�/�7�;�f���`ӯ��O�_��Lhz��L�-1�$a;���̵)J��k`u��}�M��BQm!	�����!	����9�!;��@���;;O	�<��r6l�yy�r*]} v:n� �{=�N���&��R�_��3��0�.�� �t .���1)��LNQ/��)Fи�*�4�
tt"�3��1;�E؉��-hc��+�}0�p�!�}p�#H�p��F�@���ĺ�7��a\�ə�Zf�2]���;aV�pO�qye�yI�v����d]�e���սX]p;e�nPk6�Pdg���5��8�-Ӫ��_K�Od~�l�b��i���s������Lr]�5�Qy�~�B�'����{6�f�۬+#��c�aD�y�>�4�ɹ��R!d��9}m�Ղ���Ъ��/t7���;j:����"�~f�B0�:�T�i�X�N	+�O;> rI��7��y� "'��=S� ��o4����"o�0�Wj��~(E֗4�WAu��o
�=rL�K���}X?�>�	�z��X?B�;�_� ��A��9/��qC�~~eZ�W6�b��m
<��*�)��epm��U��4���Syh��G��$FHa��Eo�V����=Z�lA���n#��`��[S�2L4<����/��(���U)�)�^ES1���p�F�y��� ��q�M��z]�La��}�)dx����U!���W;����hYW!�����2\����o/.K��YW���q�����'}�S�	���D�zƶ��m�0G�u�RS�j��9��Np�2rE�]���x9`7œ����lYb����EJ��y
OG�Nf�7�U<�� �Κ)�'�������ܟ-�/7�ˬY�:*2����={\*��r�UۜC���Z�����Nؓt)��j�l�~�g�ݏ��[��w�H ��#��W���w�o��p���p2�x[��&:/��3Ң ���ɸ�+�r��ms�k�}���e�����6~��p-ą�C:�	�ac����1����t�"Z�ԀU7�kB��a�S7m�/�Mi>��u
�}.f��/1�o��>8��0��.:�)��պ��O%�L˛��S�1�ڇJx�3�"�����Q��Κ�5��4����T���_9�rΒ��'U�9���#�߄���8Փ)��,O=a�1N�n�O��P��$�@A��f��\tbkQ�1-J�:@4`0b@��e�\���1���g��A�J�҂9�o�X1�3�QB��X뜧l���alE���4���+7�a�����^�á�ł{���h�5��6�����Y���#��vr�z���k�����TR����>�kqn3�/��6I{`ScKY6;m���ik���c�T��P�M�X����񒗚6:��'�������F�$w�p�'svF�}`b�m<�#�?�Yjn��PB��{e�T�wB�Iy��h�	���ڭ"��$)����ѩc����T�4�I$��7��9S�˸w�^|��ӟ�r8�A�Oq�ee��pv�Q?��I}$3`jʮ'}x���*����Ϋ�O�������;:��tٟ��~��6�T#J�bPnȴ4c��JZ��0M��[+��VϢB֍T�p߃sJ]����
�N�Qx���6dA���Ms��^�3����.�IQ�g�a#9��~哔^�/NW}�]O��C�ĸ;����>����<�~�B���V�W;���;�����2�zB��T�}"���TjOb��g���F��Y�r���i~�/0�aה�o �/58K��\�*-CW��hS4��𙌊�ѵ�?��I��Z��D��T�P"+�Q5!�u��"����v����[���ON�:��a�)�w##���38��o�p ���.M�@���%J2\8�P?W�<��,1������N�g�9�5�"�`���wt�9�fV���a�X�P���R�̕�� 1`mĿ�w�⥧�f�w��s�X�<3+�2{�~����:i��yg�jQ�q�%�c2�\Sݾǔ��j���Y�'���U�O륷q��_c��"�xL-q�(|� �LYN)m%A��ӥ<�]�?@��{�+��evI���N�-��p�#"��x�E��Q���ʑ����H��+o��%S�0C+8�n����l��17�v9�K��/+�Ǡ��kH��6O\~v5��4d����QK���6�$��b���O�	DQ���#�,�,oG��� l���m|���+��T	���@Ԗ��j"U�TM��=�J�e-5��7H_x�A�G���w!|]Y�?4Ұ���)nr%����wS�2�F�MM��N�LQf�F����������������>�j>$������˒��s��z���W���d��s��6g�;Z��h.Ai�&9���r�md~{U�W����w�k%-�v�p8h
�Tۀ���A^�h!��7#�c`=���8⏄��~������%�&J{�6�g�DZ�q�_k�Tz9�ݯ��W����b�"��K7�l��¶�W��@@�r&�U����+�cM�����U0P_	Z�-���cT�u���%�{V��H�<�ug������ze^�,����̦eh��R�#���'�G�;��z�v�g/��0�ﶷ0�!�i،��a@�<�C��⢐�OA0ȧbZʵX��d�R�m�X<���cD9������>߄eT1y�2-�2�	Q Lg&uC���
V�^�JǬݤ���Tv\Dh<-����C�	�޶��IGD�TT�%Dsn��p�B�v�Z�KŨBk(��R�5G�CI��m�R�S �1>T,H�b�Ŭ�����nǛD�s~9ܿwP�I�n�ɀp���'0�y	��&�s� -�K
 %>�V�R6�e�8���z�0q��3��~��Xd�H���h*�� P�P^�q<nV���-[�qE��.z�l��6T��7v��.��0����p���y�W
.B�6�8o%Y�*���5s��(�4�$b����r�凍��d���=͈տ��^�lO�UP@�?3�Vλ8Djy���EH�j��\�o�$X7�����_�|��5X���y���/�G����
�+���h��^w�gl�����=��zY��{J�ť���,6F;�Y�
J;;���
��>ݎp۷��&���y�Xw3w�����S߸��{����TN@��O�����/O\��<ʅ{���^�2�S��:Y��?M|y�!���p�-v������)��E*N��ӻ:�-�THy�&�@�2�AK��,X8^?���*З0)|~�4y@���Ҩ�XiI�VBkՉ�T"�R��`V�����.��:-C�(
2�U��&Q`Eo�l��?���π����Un�rؽW�.l��Xq����V��W�^K�6�Q���:��''4Oď�2Mm[�	O�@�aB���й�s����Qdզ��㬔1#�$���}@����(�WB$8�ͬ)��i���G(��d�8ƍ{~Vƹ��Q��>�/�nQ>�i�_7GF�U�L�7��2���jZ$ �yT۶�'d�^o�ì�7J�&q�!�MA}��<Y�r��1h�c)�� �~lcCm�7�mK�ϑ�Z�&��c��lS���V�*ϨL�x���Ň��c�U��=�)�ĞՃpt9�;�2�Ř���\c���/�.��Ci�ۓݍ��a~�u4����0Czx"x�T��)W�P��xdZ�Sٜ�;�fMS�zw�"���@8��7�~>8��-<ڬK$�i�X6�s��a��-�Evr�����ϖ���\DO4ޠBx�{�<DIdep�s�)��~���v�"��~7�h�#��&�f�$�&��z�������u��-��Ө��ITd�x]�:¶{y���'>�tM�y<���5��0����3��w����/�<��=)v$3��F�9�l��y��b��;�q��v�[C���~:�g����`� D�ǲK�
Э_yng����5?�ۚ��.�#��<N<�؃��,���Z���qń�6�
��j0���48v|Ѳ8���Z�V�oxaR!^��O�"6���| �bZ3���{�$*Lc6��E؃R��n~�DͰ8'2��2SN��f��ʍ5��!�ݞ`HA���|
�����W8⎓o�e�J��.�id+3f��a��H�do���\�;ɝο0E��޽s��K0�3[��܌a�Ñ�@��>E�:T ��^I��y-�N;�6����7=��~ ��	��9B87ц��.�l�/�����,w���s8��=J����D�d��� �J�:�0���9�N���sn6��4ȉ������4�Z��) �Qf4e�C��i|0d���E�x���ŋO%x���*���/dJ�E:/c/W�A��r�ø�P{�ik�D���<��K�[q�6�h2 _�R��t�b'�{q^� ]��C�<+�@X/ZQ\R���luc�?%
���t�ԭj�CvTmH��&%�G􎨤��[��QO�n�2�2��W�RG�~��{S9X���<�uA��9d7QDl�'�Cb88{��%�uvl���kC8�
�z�p��!:%��mư��,���P!�_W�Ҧ#��s	���-���'S�)�r|b�Q���'RH�1�եX�u�g����9�G4��@[�=l�����L�����{ƌS
��P�Z [���U�Z�T�+�L��BKBh7�q%�� �T�0���+��D\V,u�c�Q/��+�р��u� ���$���9�l�w#�n�N��*9�
I�$�N!�M=��������ב�ET��'����@I��2ҕ,z\&�C�A��o��#�lC^�$����{T��~YCP)�Y����n�����5\��I�������p��U8�E������%�y�}W�8�BP]��}&&�XE�<Om�x;}s��\�.�����j*��9>���
����J�9�6��R�$fs9,��h�U�!(^7c8�}�/`2�H��O+�K�꿏$4B�d
B#ab� ۩�%Q�.(�K� ��7��ل/2�!g"�~���9�2�X��C:�C*���RøO{s	�E��W�!>��Y:G�8�jL���.ߨ�	Y`Wlb��V<i�J)����VS�C���)�d@B�%�e��2*!�ئ�P�ߤ���{%��4�?8!^����s�͛�y��.�lӌ�G���C!��^�!�p�6�m5��HK�H����dk3#�m<��S��P����k@�4ņ���t�=�����Q{�p0� ��؊��D �Pq�b%(X��:	긲�T�l�	��U��jj!%�i�v��c�AHC���3J�)��:/GFs�Y����z�|�N�V���������ޏ�o���rZT�P�Ԥv��M����#Ǿ�J��m!ݽ�z5qi���N}�`��.�ovò���Rë�r�q��@d�%��;ry��n�����l��X?�6*�[]��~q��44G�����b����Jm����)���3��c��M��ֈb�d��J|R��X6�	E��k���iu]G���٣>QC�ĸX���@j�_1�9��G���:XD�?V�L�YB�ǿŢp��{�(GcB~�������`4X([I��I�bXGBX��O��A���t:��8ȋ���ǯx�5)�DU��W8CHbqƧ��<�R3�Z�+dL�?��:���#�2χ����)���2�}nx�d��2��Ǵ��!N���vG��t3D=K��ޜ� B�Q�c���H�̈́ $�hH5b	݁.��9Oio#�p�gx����sz�8�"W�-��c���K�W� ya\���?�D�	w�����^E'�uS��>�^M��@�n��l&�,YwS���-�0��`�<�`���A��(�6�К��p�V��п���`�G6�a��/�������?3��3��Ձ�s`�w܎��Y'��#"��<f����ȗa�y������n۷61��A|@��h�D:�����%��'�Ճ�L��z�B[�J�Cy��w���"�g�[��g�N�<�)��[5��+�u`s��{�	��f ���a��Q�BS/��P�Jj0t_��~�5
������#aPI�����a�cl��e*X�7{5��'��\�`�¡��>Oڂa|�:��)Mk�M+�n��J�R���_8�� G*⫃W}�qW���J�,\�1�X�)l��P$�l� ]a0�p\D�EH�Ͳ�ӗ�ڼe��r�v�ᆂ�Ey�J��e�
U���]Bp�����n�k�D�\��N<��(�)��GۄV3K�k3`Ut�6uur���	>}����*JF������:�����9���0��|���hd�#�r�)��*���h��{��uu�w��jb���ӕ�7��$pǢ�����&��O���v&S������ř�%�S��E�u���H�L�g+�(Y�ZH=x3�1N_/����Xd��v���s�B�ݗBtE;H�����C�2x�i%�$9��yA������|��ݸ�tt��N�n�&�T��t���A�Mf�o��h�"� ��z)�[@4�C��Y|�����{��Qa�2��nkg]Z��#;5�)��-��
ٙZO>����Z�l� �-�\�`dG�r������a�vk�nz����U�`ؑ <]I��!ǜ���ͪ�<J!�^�K��)�Uf9�4�to��� <�Z���sRÈZH���+�l�� w2�C�d���T:ܨ���C�D]|���6N��W�g!V�B�߇#�B�V��."�1��/J��7��<���F��as��gS�3@ w}��2j��!M���K��d�'��4�W*�Ӱ������O��:¶����0�����w�>�X�-�)b��|B���e�Rz)th�~A���m�1]O��5	��ڠ�0GΞ�A�#�e ��XW�gYBR8�x�jz	{6W���=�����H���B鐣�L���Y�T�d��a�r�Q�q���@�K]���a��:������/%�����y�}�a$���st�_��ٰ~�+!dut���gAf�������'�X4��R��G��2!��uO,2վپQ��[Ỹ~q��!�],�m������(Xri�Qb#/�;nP.��%�V��L����>˘Q`��w9Cbe]IA6�p���ARr�|d�1#dɋ�j��@����>���+�EO�c�;O_O�����/�T�nk�Oo�� �UATF$w�JC�X�Zn]��-W|Z���vM�ɏ�'��*�DE�3  ��+�hm���@حW���@cni`��=��栔`�
���>1:���Ӝ6 0Q%���8��<}_��]��6�3{����g���:��_˗�ew�`MO�
���Ì�����FJ��3I؃	�-�_�����%s���mչ�"�PFG�S���=
�6%4����+��� ��ވx��Z"0:�7c2�ڀm�r�߹����#�(�UP+�l1�.�������O����5�^�}r/"�!B����؊y��-Տ~����O'��t���x���p�F�,g�dj|�<?���WJ�i�M�8z�p����7����$���:m�e�O��dx�'�W�Qf��j��jg�IU���x�tjA��v^,1�`���v-oR��h/��{��1L$+�J>��Yb
z]b�E�d{�q$�X��E����<��,:0�X]7$��� ���(p�Z��-h�
輸�sϵ�Z�Q׺R4��=$N�rW�HC��N��X�M���/\��4�^O+-ے�H/�( �/�M��NT��Ib(i�ڴ(b��l���?�u�l�i��TQ��,�*g���/�i��p�0������H#�'�e\₍�Ʌ�]HD���M6�~�|;NY^�������=+�����Z͖!������-���3]ٍj,g�Æu���&Kt�r:FQt�̩�ߪi?xi.P�q�ቩ��.a���ݹKA�\���u� QRI�Ƀ�\$��W��bն�Y������n��&�O�w����#b�������r�CB��d{������M���F��bD���T_E/|�_;�G_���X�`��P��#l��$X1
���1�[��~�=��-��=`��^pHW�����9|���G��%�[���01����:Z���/�N�X�P�P������2��cjꚟ)�����B�Ȁ*7(˳���q�za^�RO�B� F	+^ )��/�)�&�>pL��|����}ژ�4)-����C������c���Nظ��M���@����k�I8����J��cϑ���3	�*��Os��ap��P��|o8 ��\��T�b��Vd�M�ܑ��ӰT��r8�K�}�0�`J ݖ���ߺ�ݖ��`�q���8b6��d�_ٮXz���fG6<���[H��M� Y}l,��߰ʄ����!���Ch��<��Њ����.Hj�ESa���L��1�)F�b�4m������۳�Ō:�~�"J�Iu��e3��"梌[P"���J�$������쭃�*ʸE�n�Rܒw~Z�/Ь'Z>Բ~�)܏hfH?�m���W#7���;�=���Ho��]UZ�����-'�Y`���FK"\v�1��W�j'2qwbDP��*�Gc1���h'���(B	8]��Z��}��$�@l/��;i�#u&}JZ�^�o�^Kt�q�Q��a�a��'fL����TT�����3���P��� z�([T�>_��\�{�Q��m�ٸ�����as�u]T�X�+�3 1�^i�Y�k\\q2�h�Ծ�!�n?�����H��:q��J�5��u+��0�f����}~���l�;{m.
���:�{��%��ֿȏ{�i��}���<6����De;�"�ע�0�धw��z�2�~�p�h�]M2�%�E��9�O�����S{��L����7�C
V���(v4���1N��숿�)REx]�g#A��u��+�
�0"Іˎ�1���C(M��įxZ�s=�q�Dw��?�u����%Έ�l�6�P?���@��_CD&vu�_�~U������Z]�T:��<�9Ry� 6��Hj��RY���_���95?������An�D.�q�p5�K ȣ�ƛ���ئ��sJ�@W�"Xk����9[a��'��<�C-q$�4,WqBx���o�u$
�B�(�s��b�3c:�Ѡ3#N��#L��*Y�L��`��l�A��f0lH���y���ҋB�+\��߉��Ud8�Q.�b���қ�@Z��I�h-�^-nb�j����V�,�&���C���R1�a�4�D�ȀK��O�j���?�W�Dn��O�67	�R����	Jʗ�:-�hz�S1���N�s�<;�/)�6�
eo��؍��,��`��N��{h�޴�����h�v��TV�~_��A��H�rAE,-׶���#�Y�����ǳ#�6�t$�EWXV>G�(X3��zZ������Ԛ��D#�A!%�s'�q0` @�P�T�[f��<�h�ow՞0%���Q(�f�t�R���Qm<�J=��U��V_|:�z��8Z�r����K��`Ğpy�=������oj��Yi{�/�0�T��3V��m��[m�������K��8��7k�Ei�@�ɏ�
φ���Ra.�G�r��,R-�.s!�tЍ1�ݸ��*�iP�5����Lt�>�����K���y���V[�K�A!M�?��N3�x}�k�f�s�v�ba@]����_�65m�j���! �����{�b=��cW��(aΙ���C�2���� ["���&��d��)+�(��{!�Y�� {�5�V��q�U�E�ۗ�J���5;���ʇ��N��J��a�b#~Lٵ�i�j/�p�Q�R9�j�"|
�D�9�t�7���ޗ�57RX �x���b��*���ҵn} �hh^o������& 92G�[�ڳ��NK��F�����C��3z�<塮NY%��<i�.�̃S]	w�<�L-$R�=�t�'j?�mY���]`;���ߞ�O��0���8�Ǵ���e���DG������'y�FMc��pe������w�l3�NT�Rㇾ���Y?,���,�/�S�k�ҽE}Q�}wyj�r���c��e��0}^�;��"��%�5D�3�O3�nL�C�i���rV�4<�`6%�ǹ��xx�B'gs[�2��g�Ї������!H͓:�� (�茦Z[\ ���>�C'���T�_����A"�;QMb���=���kE��=(w��7V?�����<�q�̖�'I��-��Mt]8Zm�����l�O�b���gV](�J} 7�X%�L%���xZF\"})�Pqtf��k����c��8�HT�[(t9揌 UB�*�7�����l�r	qί҇�#O��H�  ��^�hKa���0�~�^�|��y��m�&8-ӯ���W	��k<`~%k}�r�E˒Y?��v����*.�= 6AQ�Gs|����xn�i�@ E)Ս�����A� �N�9`�1.���D�e] �[�{�$������1�,���߾,hD���Ҭ��c��1B�`P��Z���;6>!*�QC�i��.p=� ��e�2��'֧�i!�T^��ۤ�����0ErP��"�L|�t7�85�)�w @7>�aVV�<vɅg<~lo�@��:�b+��r�?��5 �N�8M4A�25�I��I��s�%+Bׯ*�#�L����~V��GoCppE|��4����/�UvB=���<�j�����ِ��2���1������8�W�,%E�1���n��^��a�a�ō UA���V}�Y5r�
Po�Ҳ�����& ���#0ۭK�ԀP�.7�eާ�*�(�~>f
Z�j����Rpܡ��!g�﹵�ߝ1�y��_Қ�.�EBO�&Η �l�Ef/r�vYz�0Bwލk��݀<���u��ҾHx�e�]���K3R� L�f.o�V��k�o�92�^H�9��%����F\�?�ѿ44,�8Z�y\�-�$1�:W��R���jd")���G~��������~��i�r�X��\��c���Ʒ�Q���=�~S��ǌl,:���i���=Q?K�� ��?�@����׽ojI��"��Q�?�ק��E2	Än�=sgy��W�l�C�0�l��N�6O=�]y�f~�K��UVh��,�Ջ����%���fn�2�a��靂%봥��җ�7ZtA�N��,����hGMLQ����0
U�Ϡ�c��'i�cbyIw#\=�`V~N�5�������	��J�k����Ь��Y$0�~�s���%ͮ񢅈��%+z�F�i���8�2���Zքb�����5�D���3��n���q� �v�64.'�
�"��đ�}�ᓋ2�epx������P��%�n���-����A^!�k�
UU����Ѓ�d�j2[e��V��d��A��rdG�-U�l�S�{��-�v�,N��2v&"���O�9f�SI>��"�y���<��f��A7�N�*X>!�Jc��Hv��VRe���SA�R�.5�%x�^�k֭��dw%�T�n��Y!LN=	Ŕ�g�b��CH�}���ǃNA����=b-��ʠ���'���W�=�V0������e��{=��(Y�1\��a�!��;�YX�� ���?�)'��	�0`��t�g�t��Ncb����v�~��W��\���d��<��
8k3�;��|{�W:�i52����xipy�bק�;�咑�)�U�5�x�7�ֱ�U�����t��pNX1ǵ���Fm�2K��s�݄[W77du�U7n��M@�-}Ǌ�u޼��+�d%�s	��I�#,�]PB�z����ma�:-<�:3P��1��J!�v2?d�v9�"n !4���*$����]	!�����+�Cc��E�~5&�e�]�]��s�_F9#*sH{���>"�V]~��b�9= �����������YQ;ϙYD��Aڑ$ �<2	���	{]�[)ؾ�R�1�٘u��>����FT!h�*��WIV���9Dbϥ��|b���*�"���>� ��sE�xW{ �)-]�z\�t`�����I{�]=]{��q߭-ca�1����Tp�h�,G�q�P<�%���q���a��Kͤ�7��j�}��Y'�������j�"���������8E Ȃop��I㳏��Ff�4�O�����x�{�7s�����`��{���?��'��pHc��I�r x�����|��o�0��Sͻ���{q�����娐o���B��~n�dKx���D>��O��ɳ�Z�"�<��z� S~DI�Ň�x�Q���$���*��w���^>��K9^�ժ��N�쵟ɡ 0c���������j�Q�@ټ���;����ǲUS��X
q�(��Ô��7�M8y������ၴ��P�B�J�3��T�D���ޫt�[yD�V�Rh�|:�JLԬ��^��Q3��|�4O(�D��Y�[�;� ?��3Jْ�{#���P��C���d�M�i��N�{���_}	c�(�K��W&Vs��qMg�T0��}.sZ�I�Dr��"1�4��&��X�C~PXQ���/�5\<_�����;3��i�q�Mh�5,ȅH6�1��~����*g/Fx�	ף�ĎJf�w⹳T���өew#��҇��vGW?����:���=��Rw��[$c_ߗ$M9a(/����ΌX�yP�u�z�3�N=]�n䔙Q���.��Q�CV��&�=�P��?��oz�Hj�����H$*��jH�`��?�׌����������ݵ�S����i(lwb/�7<t@�~,�P?���͚A�����Y���j�*5s���S=^�%���{���$�^��NL�ې�ks�a��*���}�
$�qe�pjA�m�bz�[<��`s�,� 6�=���}��xzY����'�����d��C�
��8��<��1��s�v&��ĭs�]^�صf��s_�1e�\��󺩢�9�H�IuyZ��6�ԁ���ɡ@�~�b�1�l��ϩca�O��B�з��s�׼G��2�˶b��%�M�ێ«!AY����Ik�(�0C]��煠�)����k<�~���:�ëQޝ6��遢f?� �L��9o7���wP^E�V%�'w�w�����7�{S��C�I��k�W�R䆡8}wP��ͪ���25��~ɹ���n�fN~4ms���<�C�v%��$U8$�a�RW�C��oЛ[�4��L��ȁTaa�P�1?�Aܸ@��:D>�OGE��rI�Πb��4vW�z&�:%�%��~z<��R�!5M\~m%���
<T�L�t��-Hȳ\OK��o�����Zk��X�J7�
�{�p�;Z0q��Q�y��2�</�g5�Q!!ʳ��H��5M/20��� �n�>�PN�,�0 G�l��/����*$Z��!����<�k���#���Bb�v�YAu� �|�P��Q��s-�#�����R��P'w_5TR	1�uw�6�BÁ@ �-�[��6o,�����_�P����2g���7�<�K�Swk��}�d��EW=�T_/|?�%X����6�.!"o?����'N�e��� �H�~,^�>�� P%9ޞ�V�S��g/KWn�{E��������Wц
�Nݶ�rv8��񞨐<#ù �E��G�},0����BA����h���#IS�������f�Lj<r�F_�'�M�~�#ƨhJ��j��#���5�O87E��~yT��~�S��/q�@�rƧ�sp���G�Y��I�V O��f�Bԏ-n?�\m��a(l/T\
r�0�ֱ�.x�z����.=$(��o�g�Y�tD6�ӗ=vf {7)�b��fDUm��Z�!G�.)؂��o:���\�[�!;H�~�h�4�ڒމb^�Ȩe�{8t�O� �>(��\ağ�ү�E���1&&�SRE�]Q�5�l��i��Vy�����o��|�T���P���g��x�x�������E�
�e�9��}��`l���F|�J0�A�w��k�ֆւ.3<L��"#�]WLN��>��<�!ͅW	k�E�6�l�+�S��.0���v$���MK�-Rߩi#خ�:���ߦ���8��q�NJ�� ԍ�Bc��������Y��~�8��¯h��ne�ut*�����*��p4;��1V��d���j��RC��`�����6�$�u���*�1��uH��i�凰1;Օ<���g��V���g�w�]����n�c�Lz��]�N�N�m�8�R�-J��8
i�iÒs���[xϮޅ�_P�s΋k�o�DU�Uٍ.1�-[��,�ҁ��L@�Q��7�P���,14@���3�Z�Wd�4���'сq����S��TT��d����=p�K��Q��W���n��D��rJ����`�i0��q+��4$W�� c���d,����B�ԯ�^�$�.�3<�|�c������LЉ$����Ĩ)���,7c�uo�`�7����=6�c�s͐�����������+,g�_ϋ�v��&$�H
=C��6g��I�Q�<�=�Y"\��ru�j�%<q��#.�D�B0O����'��őy����݉6$�6�vk��O���Д�,�z��4�D�S	��\��y0 pAC�ŵ$F@�s�j�3/Zx�����;8����e�5q�,�������jB��#���ra.6}nQQ���re��盞�t�k9f��Ou�����<� �M�o�B��<��J�;Վ�7��������V�Y��k���>���R:yH��y�(��DhmSkjh+B��dS�7���x��do.�Y4�q�A"ۯ̹��p�U������#�	՗����%��[���I��k'��FlfƏ~�,��������R>����0���h?�쿑�6�����	�h�"�m�_ Iϲy��b@w�߷7����ʬ@�b��@�EFˁ�V\�C�kҽq����x�pfo��Ś�p��P��Pia�ѦxGG�|Y/F�T�u=^�{�Cc��+N��&�$0_�����FM�=L)�;�ޖ@@�M���C�������(��u�ĕ��%{y��0�=p�~-�wP����y���ű4�}��q������Ζt�����s.��!zK�d,�K�M�8_ǘiD��xkN9������튘/r˔cV�j����u�W�T�J�߈k�t*jo��f���D�-��t\��n�����03A���9�.\��wx�������xQd"��qM@^%D�ˉŻ
���n�c�o�I]��i?��П�"H"�s�(�q��wǬ�zZ`Ń�v0�8�������@����4�5��~�ޗ��Έ_�=`Y-Az?|k� 0������C���J�?�!�u��;6k��z��*�5��4-��f0�,�g�<�\��s�q����E���+Z?�/����@GG����\��׊�J.�1��!W9zv�z��O�#��c��+_���Y�	W#��S�gc�P�DF�a���\	N���%V�q/�yX�M���?�W���-���L�~8��|qt��C�T���[��Ro����`?ZkL���WPCe%���}�,�ɵBb�c��Tn���g�!{�U|�߃pM|Р_j(e�v���JU��?'�2����i��<a��Rm���R����i��ڃ��!ӱ��	�e̔G������8�)�7��4]*p��Hr.�}KƷ7?�'<���*�������k=Go[��&"��諔t(H�W���Al��z��Ya��ߗֻ�����G;��*߅$GR��H�-�d��gH�dn���E����\����)3��Ixt��0��۬ ��越M␉mDV�I��u�"���f�
jnE��92�B����Ca=C�!ʒH��<�X�'�����"2on���&Uz�|��\m���)3���n�۲|BS�EO�h�����9�Sɿ�����x�G6���.�	4p���؛̂"�����?�����N@q�8۶��zH��`���� nT3�ln=r�q�7M�t���%��Pmi.IJ9$���qo�'�m��v�]S �+�7�lQ���|Һ��H�	�9���w���)A*��2�9%7 �SO���t�'�� ]��tM$I�-�nS��(G_C$?�7���]Y\�ϸ5Ғ��� �԰��|���lSՎ�E=�����ch�`I�9��[�q����~��&a^�/��anF�1�H��S鋳W��F�Q'�Ֆ1>��
�Œ�]x�;��`��p�i,v�b<�$+��JӏhL��͘��/zd#V�����e�	[����u�('�*�ˈ�]o���_A�r�ҖQa�!�r�1��� �JG;ol��	c��]�;���.]�~�E�"�@ )�R�fbc!�'��|�%r��L���!-���5�P��O�@�܈��H
�z~��&-��Ȏ\O�U��鮞[��"DOmS��п!W�!l~
�<g�S3�ܻF���ӆ���(�%xPF?��C���C���{g��I���`i[?u��Q�%�k<�wZ�7[-�bf1 >g����g�C`0Y!Юt.>��_p!iY7�%9D�é?LDe`�� �fY7ıg�ҶiO�pJ�WarS�Y|jdq/����C�^�unu����9K�I���׈�?Z&X|ˑ�&��-��&�]���Gm�OGw�TԜ�Z'9��t��V
sꝕp��|:N�)i����v7�S�6y�[�}ud��W�	^^����з��D �$쐌�~z�wS��	?M�s3��ds[X{�7gLU\�l)�јm;��\W /��Z�7������ϑ��x�˂le������M���ld�Dc�҆������>4BP�8øiyM�lJ�,6Wa�y�?��{E!�n�&7e��ǅ��oi������=�F���!����ɝ�H�5�S16�K�:(��B��Ƃ?��d����V�&�^�2\e����De�������	�������c�ù�0���JJ/��+�( ,���%�j'EL���%�A �'Pr�;��rb�:G�{�ϻF"��a�|�-W'��r���A3��yJ�ju��v������K�nE���o��p,FьZ)�tV��h�.(���c��3��K�9'�a���q����ֶ,�W�9�����\w�%�!��ؙJ�p@6dOѢ1)�*)�PZ2G�N��1,���Wb�v8a�����	Y�@���g�qx!����΀�X�t�`�·�tx�Vu��*E�Y?>��y����"����r!7���8P�]>����@d'���WV���:�M
�Rj��`a�����@���"��5�~֒�}�ë���@���&	*�m��6Y
cK2�X�(�l���3���}6S}�3�q�>̣��:<v��f҂��=(*9��g�����﹜ytt�b��v������9`5��Rys���lB��yȌ�b�J�,dӪ�3j����̫�9?c� l����\�dL-ul_���~3V�P���*o���ńi���]�~��[�gE��O���i�r� iC 1�HQ��߽�b�/7q}�����
���*�:榡{�����i/�>䃚�e*gָ����&R+���1��c�����LFT8��DY&�Q��y J�] �^��p�A��>�}L��.*�#�w� �S����+��?D�7�4��O��	���7��{����e�Dt���uO+��%E8t��X����6v�̚B
I��,W��1��xyҗ��Ur["��g%X.����˚;O*�{}a<q�|:�T�n��V�-8�qgK.�TQ�.&�2���_$�c��YKB�أEp�Z�'�>Y�t��t����I�ȝ�Mn)*�`A����Z�ɨ8>���iIs�=P�j�����X ��p�iI�X�E��Wr5�B�oZ�>ddcc�G�+ұ���s��l�h�DY��ތ�o)��a��ǽ\��&���:�����Uw�P����7oaX�[J�wO�و�ȧ/(��L��uZ�L\���5A�d,!&�aR�A�<Ϲ��':�0�����OwJݘ�,�'"��M�?}�1��n�|
 ױ�����;Z�X̓�����kz2�Y��Q%Vi�l>*��KN�WBv�ߕ�C��8��S�|����:,
�<�F��4�������d~����Z�n�6oD�-�P�6[LD2:�b녅׀x�
-A�15d�IX��S|�L=���1U��3-]ʙȏa�MĪOQ���7�Kŝ���u� (�!"���wr���*�r��ew��&�:�q�o�9?sň7Ŗaqٴ������R�1��!��!�K%/C=G�F橚�㩬Q�.7�N����4��٧�-UA�S�R��A"D�Wz�n��fd����W|��Z���ةF7H	J��Ftlibˇ&�ō��������t{�,
G)�8.@��ρ�n���8gL��'����S<��Չ(j��A��`	�O��am�1(���v#�d�*{�{��s����v>��[�L���Gi��Y��N�����܍v�K�b����s��l��iU\>whw}�u�$Q����/Ѡ���#�X{�
<���"���]s\�_���aq�R�;_E��*I�K;�A�s�>q|g�݉�#���T+O���=pو�LSГA�_����e�1�� �O�Ys�|��G�Zq�m��9��dT��}M	�M�1�7��a�'R4�|-n����G��*�����-L+�CùOΨ�W�����{"�����E������x D'��J ?��|x�{!}�I�a�mϟH�*$�8�c�5]�e`�&>e�k��6Ù��a��o�L�XL��ѱ}����8X~����N��G��.�[x��ݔ<�̿�5���o�����l�@V]i�}&����O	��d�f�Z���@�8��_�5�c�QU��t����� �3�Z^��VO렉���9�OjY�VI��6dќ��=7qJ&�1������ޑ������mPN�h=�U�N�V/��l���6�`޷{z�:骯<�	�o(�z�X�!j���/��o����~r��;ܕCr�O�}}��z ���HL$뀕�+��v����n����>	��.V��c�5ؙ���#Ⱥ������>�#�ZX8|``[�ɏv����b��3~�`#,R�x��Tc_���`j�և�t�)�W�������,�Q�2�4�H��dU����VzS�`��c�o?�:<#FZ��P�K�H8��t ��-�͇�ױlO�|N8���#�����؂�m��Kiഽw��2�{~���{uJ0o�=�^Z�j��~����-`Q�U��_-骤�i���ˡR���G=�eO$�~P2C�s���W���XJ*q�}|xR9�+#�l/�QF��L�#�s��mu��abu�a3�ٚ#�^�dfK�%`J�]T�ýJ�������T�%�3��&'`0�j[w����!�@����|=:�tlU��gvޗ|@��AV���>��7$u����=����H��TE~'%ɶ�2�>�X�{u[�Rk1p����*��F�Y�%��̢�\���<�f����@)m�O!�,0�=ΐc�@Ύ�ѣ�̣��aP�Z�a?Y�X��9���S�?����U��ǊR]�$57�4��;�c*Uk+�r��Y��;M0�t1��t���
�}˴bipl2���]�+��B]�0@��W����K֟�P���)k�Q�b1�]�V�aſo�)�u��	l�h���m�����*R�\n��̀��=@_"��gЖ0a��� ��f�눁����\����!I%{���ef�8���|%5\8c�q��ibde/�
�,���������6��]5���z�	=(�$���^ S���x��w� ���W��6f>ˈW�/�o���x���3�Y7�c�LX�о4�{n~⑵�a��q�FHR��u%�\i�Ra�����h@+h���d	l�8H�X8��_T�>��Λ�K���
<�Cʦ�t����拤¦ɤR������Zb�z���,/�Y̯�m��~�~���Ѱ�7�5��~8#;%-��I�\G�_5�̝&�ł1	��`}��yj1]�	2U�j\:a�a�%���mKn�D�{�I*@�t=���i#�צ0��鵎�R�,�ZwH<��O�Y:�˿�]�Ul4�#ތ-G���݌��ʹ!/N:Lx7Db��(��V�
��3��ާ-*gF::�t��ǜ�.y��A*fV�Y�Eg+1��BuU��+o��{,�Z,J��	v`8�>W����/�Іn/-}~�Q�Aj�Q�e@.�f.\����O�Ǝ)RZ1*Fz�+�L���𓧝����!�^�p�Ų�������~�p�E��D�Wp�����;q?�E#G"-�u�I���#�����k��l��b��p�<��e�DL� �E�4��bP����b�+~\�_f�U����$Ԅ-ʏ��,Y��;������
S��S؀����W��)�F)v^`��)�y��A糸����3�(�S�A �ԃc��
���b���;��������p��0��S�|������Н���W�fu3&��;�m=ڨ�V<�1��ӰZ�0+�~2��Z�����:n�.�g��j�[��֜1qH�d��.�����'�����_{>E���������L��+�$����%pԛ�)�-����)(�q�$`h�ga�s�KX8vzs���'Bl�f�����e�5"(Mvn+�jy;�@˲�3l:*#t3�(��� ����o��B>,0~j�W:���U��Kd>�i��Kf�3���h|�1���+A�<QlC�Z*�p.�b�8`+Q0��J0��C���E3}F�O1�\�"�X����ᅀ�LKXn�0s�ƒ���<�=leD��|��xV�b_� ��M�Q���2
ZN�G�MD��6~�^V񭀪�e�긔�j7�d
��x�$��n-�SQ�A��ȢD����K�"P���E��T�*���ֳ�H�KFPf�E*���m_y}7A��i&v��4Eę��k_6$W�ys��=����#5��zI�͊�Yp�dj6-(�pE(������a�:�wBx\�7岶X�Sk%}a_hK�t�����`����L�x�\��f8Xs����Ԥ�w��j�(��ט0+���{C�uG��U��Y��>ur�V"�����k���[����}[���b�!@�	��<$֯߳6_-<�z�( �x���ԑ���د$:�o��!B<��7(تp�?�8���8.����Bw4n�r�nuԹaP��w�~;��L�S�ȇ)|��]�tZ�v�������l���8�Z�fa�(t�l��
�8a%f���P�4��*�^�η1Sڵ��$Wq�7�_��=#ط7h�:��������I�r��'q�k�e!y����� ��� ��w)X|��wRM����W.����uX�׀/3^��\|�_�m��-��g�.Le�IGr��]���N�.�-�j��^�J�X\2ۦf�&1\�m~F���5󰝨&�ZrÛ1���䖭w���p����Gh~����D���1ŀ��P)�J2�3w��X�}TK�1J��=�7�	���ˀxQ�b�[��6 ��?&�~��*��GR�@pSQ».��T��d6�Q��.�)Y��n��I�c�B&� j��&J_1�sgl؃s��W7� ���x���бӓA�i�mn��������q�.��~� M����cϦn��$;���2���L�^��tWl����%2�*�(I�������S�A��!�������q�x�ݛ.})Uz��W.�Q�ѷ����r�Լ´�~4���y�O=��Vt%ȵ(n^b{%qfE\)� �oy�-#�Fb|��zc�/�����l��|���/\��Mז��-~��$�� WH@rX2��b!hIVLǦ��ğW�����M��� �B8J����lԌ����HtƟ5�����Ϭ7��-�=0�ٳ�E|9n�;�i�����bj�:.?#�)s7�b*�+�S[��Qv_yP懽#��`E��������o����k�pn\U�[�5��SA|�V\����v�\\BfŌT�n��u�JϢ��Q������ꄜ��*[�y�5OϮ���A��3=W�W%T�>9B�@6�� !��b���v�L3�����=s�?�r�ӥ#�C��_*�	�g_��|Qp!9!��vB���WVrĄ-���ۏ@o=���gq�g��=�a�0?h��.T)m1�"t��Mb����zS�	����^����
�Xw\v|�%>� ��� r�'N�/��	[�5����~M������\�%?��(�V�.���$���9��'WR�і�"�n�%^Ʊ��,W�w\>�/D�I�&5Iþ�4`p��&&��<��$M��������Ґ!)gh�Pʐ��}{0�d�����On�[���/��g����;�s�ZpTEg4�5���.�Nx�rD1<*���5�43?K���I��G��%b���h���Q:���~�<	��g�%bn�]�/�<���^��\b	L�!�A��p�{���T�&dR�[�FI�6���g�� �X�kTt{lD;ʆ6��VeoH?bH�v��K"&�]�<�	�B]D���b_�S5�!��am��*�������mNN���)�E���\�"|�.�����QO0�x	���#
fH4��sH4É�3�+j��t{mʙҔ�zlX5H�ʓ,���I�FW�~à�?;�]N���8d�b�;���>�Z�цe�)���7�?}P����I�0!I)o�"��q{���F_���Je�U��Vs/���$�o-ʬ�Uy0��5M�ISx������yb��Ң�B�,� '��U����L�H��P���N先�l�~FJ�a�0:����keP��E�ق"�đ#�=]��)���y��V���m���Jf�s��A��|Y��?+陚饐����<&�v	(V��e�gM2����W��<?J|Q�U#J��� ��'Sڻsv���1�*���A :��S6ϷZ�����9�z0o�tu	lg�е��+��G���J�0jQ��9�h���{5���&�S���c�O�m�f"�.\ә���S�37�+� ���+C�M&���l�]�����m7��2l3S�P��d���-�l���zA�õUei���jL�;,���	`�Q�A��jݿ�"��0�].p�ƍ��7i&<�)�BE.?�m@z�����I�>�J�߳���g�d�;;��?�Y��-�E�������)zfQ�4�D"/ˠ3�Yl�gW�����L*|�~e��0�`����MxBERZ����}-^����m�kGW7�=����<�]�'aߙ�LOd�%�Uk��R�N��@�{�5��+3#����ɹ+=9��-zp���A��� ދR��M�"�M��q��>#)Ԙt-��꣼�I�8���J̱P$,8ڷ�Ж}�,�e�@�_���kJ��^��.#E�����l8���r��o*�59����?�����F?���%]$d��	��I���Z�Ƕ"/\Z[2����#s�مq#�˞����%�Z���l�,pq���T�[�S�a��QzㄊnX �-����b'�Sױ����	��:�%+3�r5j�90F�F(d0}�lPL�𣶯?	�-�Gp��Yu�j@jĭ㪛��>6<��i��9UI������al'��,c?y��@c�v>���%�{�������E�|bZ���	�1">��(p�D��cd���j��s��9�wz���D�b�C]j��B^�'g���ߥYBN�m,K6��$�~����|u�̨���~�<� y|<�8�_D��č��z}���>Oaa"F�+U-����_)Lq}Ѩ��"��-��P�����>�m��)~!+J׌�)LfA'�AJ�}��v����C���4���]�D��Ez��TL^�L��Z����`OFwO�Y�^��2���YL�߮ZX�~�;ĂSy�CE����\웮Sc~�"�#h����V�K����}�\d܅����Z�V:���;�^2#˛��N-t��Dx�Ml��x�*��r˴V�(`+��n��!���afޥ�2㵭vz�����J�����fj�����'79�dO�sSųD�_N8�ח��
�XG��ʡ�߶�`��W�N�`m�>�v��ю�ű)�Xw|�w4ō���&�Ci�	�|$��ɪ,mT�i0�(n������`,�״�����bý���ݼ~ZX����.l��`Ð�S��Ihd��>`Yק��]i|�JG��n��΃�rK��@��������-0�R���I˯K���U���L��L����9���C�Fۿ��Jx ]�����v������� �k�5xrN<eYy�?�&���9���e#����A_/)��r&�.b��ߧ�mmw*�"��;�|�{k�7pԔb��l���T�j��փ��F��%Jq�%��;];T����HV����u��V�ɷ�=MR2ˬ?��wL�0Ħ;^Ri�{��k&U���[y�v{�^�BK�����cςrc]^/�4`_ck����j��XG�RMX�[VTw�As�1���ȸ�q���x��50������(7�m���c�!4`q�eV7�T۶�㤨��Y5��a�'߰�Rd<�~f��r�Բ
�iQ���p��&wkZ�/<��`����#5K����`�aSA�B=%64�+) �H ڦÞyNVP�=צ��0���	,'pS�	��FM�i�����.��Ǥ�lH ;��Ҥ�<��m6�:����KƩ�S:B��� ��:k�D�7B_Vܻ��*�D�k-��b�٣�1�������F]� �N�U�fI�w����25Z'y<�rJ{`�}�u�W�z�HTW��-S��R�>7��\Y:��|��`�+��Xj"\��蕒�7�������
D��FH^��h���<C�8!���<����Sw�M��Ď����=�Գ�_�_�b�"O+��zP��La
r�#���`�Ys^�=�A�^Z�b ���
��=�""3�gʻ�Z
4����[#��_����"2ӻ�#Z8l
��3N�2T����`:?��S��5���:��۫�,������r�u��!���T�x0zb~���;k�8�_��?0^1q٘�Y|T���D���SS�(r2
�# S�v��|G�����K��Y !�}'��U8aF�s~���_�'Bk7�$��ܞs����g�X?���S%o�03Gۀw��`(��󍻴D�<oC��P���1�����������陛	��(�R�v��O�Շ �7�h����Ą�4�_���C�t/�|�&�%�IO%��8^���f
����O/�Wj_tP��ގ�fg�0gf`�,�*N�������{h-+>��a��9o�?Q����ST|F���Rvz�r~�]���n~Zȹ0t�t�U8��kޖ~]087r�-�Π���g�����O�9 (�(�/R3�
�� PT�)C��#�M��l+}A�T?�U���g� ��V�W�����T.잩d��^��D���.�B���;E�S�JeN�����JCkD�{�U��oD�6��%ޘ� 1:��W�
�w}���?e��(%?�!u�vד>������~�ɓ@�Ȩ�ʅ�r����rXh��y�����xs�d�����q�`���بВg�a��I�dۊsb�"^u�J-,x��x�j�`��r�m5����Q��2�y���
M��_l�~,�����H�~��=aa�4����cOd~_X�N���]�K�]��M��>��0�>6C��s�!�ۻ~���7_I�ό��Z!l�q>��T�DS��;��e� MNk!C�#a�Oo�{H��a�cR��Sj���G�M��}s!�ui�;it�D9Lmx�DH)�}!r���f7��3�`���sslPT�c`ܮ%��ϵ��)V���"���P�RL)�l᝴Q�Ɔ�W�5�@����'w8n���֥�qO�w����Z�_���d��ۚ[1{kb����3�^��ܿ����N
���=�ǜ����*g��]��F�m��OAJp�q��z���.���	��ME˷�:	�p|��K0�n����
��
�ڤ�c�%nv#���B�*
����M��X�|��N�rF����!P*Y�H}X��E�d;�"hp���a�[!򵤼O�l7M<����AE����N��k�b]}Z)-�<G��~����Ozy� ��QH�R���R����]�%�h�S�_^,χ�!�$���&)]�I�%��;�������́�s�J���)4*�
0�X#\�BƓ�[������1!F�|:M�p��N�CJ��X��
܄9D[��s��N蟒?Z4HB��}�%��9k�F1ѿ������;z�V����	X���l�oB���e>U�|��	��EyC|�k�NY��ɴI�B��a��	)�8��~B�m���G��%�jrx����U��3JG;�<*6�w/E��5~�� ��} u� �p#E�#�|�s�^�X��� �>{J> k%��M��UG��jH�`�g�@���]&��Db��q�A���5Qn�ĕ�x��;��!86��!�� �YFk Z=;���U���n��!���m���J�W���hC��Y&w�eb�������h`(s ���ް�,Ub-�+�EUn!OYi�P�ٌZx��cR�ʼ�>ݱx�z5�|"c/fnC���
������"h�4���l�W�Nd��wV��k���|�S�J�o
ᱝ���r1�b���=��=��~�f��nSW鵄S�]��o9:��+)O;"ʹ�g���(��R@��DD�e����ҍ� `�JQ���u@7���3?e]&��bQI�&Y�{�D)�	�X:PL�{�XE�q��d=�"ї2>��~��x̕Z�~yih!�Pf +$3�6n�j��5���Z��Y�6�f��a�/�|�/I����By��੠ ��ذdb�Ї��?��VK+�ğ�� �B�ؾ�=�L���>֬�gC�n��g��KeE�7�P��˄�P�W�P,{�|��CQ,cg�ˏ:��
�]k+Kp�E�4ꦓ&��}�0��FyW{�_����M:A���;���K�T<`�3n��}N7�5'�Ǔv��]�6|0�/!���f��Җ/�:i}��n#�����ǽ�˅��>��=�T7~���vbb�+��n�w_ɂ0WAx5/�=5����,��(S�`D�� 
tZ��"�u�~�Y\I��|n������H���s0)I'��RPX�"W���&��sk�{[_��K�i.({U�#�����t�C*�����Ce��b�}�T:��p�_�����v�;Y�5alt�,k@A��	6
p�
�x�rd~\�.Px�{���(�KDόRe,�Һ�z�h�����0i�#��_UtX�bh�wG#���j��,3a��q�`g��O���&X~Shl������e>t�ߕA�݈^�[�`�1|�$ڙ"��ϬЅc�:.K���̒�����a��1��q�˳?�hJ�^�`V���`���Ge��.m����\*^(���kͥ��e	� ��U��Fb�b!b�|��V̖��@$�"���7 ^���Z%��Xӂ���U�=���;�"��wf��͓҃�fI������*�8��y֦�M0X#�s�"%�����ܑ�0�&NK}_lZ~�ְS�I��C�p����ږ%~�/����	j[�(9hR��F�&�1�`IG�Y�j������2z~F~���@��n�0a&����D���q����2����3�Ŷ�M�#'�A\���}�2�M��k!�|�fyCX���ؠ�f��+Q;��F��ұv����c��yՔ�x�Ϯ�6$������}K�Y�7~J���1u�35�or6����!/�������D溗�h��r�ڗ��Y�c�i��*"U���{Ra����~�%Jcf�4+w���L���E�ѱ���p6�A{���'@�@y�OC����2x嘶�[�&G&�4��i���-�Ƹ�T��6�b��'��xg6�[��[۫��W�3�����pt�-6��e;ec�K�X,��D��3`��|���9�D �%���6�ƴ�rG���8�G�4�@W�?%����%ukU�6\�m�!��v�`fb�G�I+���q�����&�*H�����	�z�}c�j�uT[iV���?P<q3��RE2�p�|l�@~1X��b6O����ZtE�����!Q6�M�Z��Ī1V�8�c����(l]�8���ߍ�� �o��Q��ɣ7d���@�S�hz�Ҡ(&TaOS؝��YwM�m�Q1�a�)j�l����1�q;l5��5 P۞��#E�F���� �ݤ�4���2 +D4���^1��Y)�@���\�Mp�8�9ѧ}Iq�Ab£)d��0X��`L���ڞ~��8���˘��v���a���y����s|�=nBΑ2�� ���F����Y��U��ȋl0"��Z��1�_\���0�S,ipw �\I�.|r�2����[�]��K��Zx����U뭂��� ;^l��A-�Ǽ��k?�8��^�����ejK��K<�!!xYKu��N�0m�p���˪B���^��2�f�}�Vn�Xx^�� �F������V��ǜ�/�#���
'dj�O�E 棉�`3TIu𪋎;&w�.I�.�{�r��,1��G��ٝ���ox�����N�xc��s����Y5Hn�ȓ�i}C6e���l�}O���'!��_NuX��s���&W�Р\<���K���2�'�_D!=��ZI��ս[����S=i9#�;˧"�d
�ie�03���T91�5�-5~�I'���Vf]I,0b�J��p��kD�R�O��dO���IL�N϶N�n�;�R��R�o�"��������.�?,5��l�:6���V��qֈ��Q[74��%�|�Ё΅I�8� ��#ڀ��n{"�?�����'Ry�:�J"�Tu_p�B��HȈӠ�M�6^�vL���ߓT�1&�8��u��=W��?ڗ(������	�?�W����hc�rL��;,�U�eoM�k����Y:DU��ࡱ8�Q��!�oYĤ�v�QC���L&0%���#q����;:Gi�mX�������xwR���.��g9���1}��Kh$��0Z�l`� 3���p��z\��iG��������eH��i�6)`;|����ӹ�D�ֻ�T��1��<�;���f�c��B�ռ�7��Oʓ�iТ�:�c��.��!'�B�øn˯�(���P�5
M �P(���Uأ��1�o�,+Մ����T�|*���2̶�.����-�wcF���덛B�Vx�ITܓ2V����0��]�N����~6�����<c4(���p<�����2$�����Č_Z���Aɖ�#Ïq���e$'�S��n��Μ�$N�s#?���u_�CM��ح��;"�g��n�ƥ?�4���OO�����"��f��|Ő���C����%,Z�q�L�F�'_bK��g�;] 6L�"��t'aʫ�9��Uw�b�h�e�&ץ:k�ۏ�$YYu,�j#�v�)^����uӺ/�_����(��~W�cene�W�f��Ml�(�>`�*W���"'{q}q�K���aV@qh1��z�����	JxC�a5��;tg>��Y#��5P6�A��s�_A�����Z�+p���	5�b��q����s���s�>c	l�a@y�Sɬ�'F��Ƴj%Аݱ��:��@e�d�����ͯ~��MA�����c6%%�ȹw%���#~� �ߌ�]C��<&#p�����;��=�SV�xd~G�o���b�7�_b�Z�i�I��i9��Ѵ�|�:5KGwMv'��X�~���I�KkP7�\�m���J�e����#�����H̛&�x>Β�k���X}��|�|�P�`�j�P8��a��:�tt���x��"`j֗���O	2a�ueo�'k�1�J{vV�[��8!����ww�Ty�������s����4Zw(����6ZL�W����"�����j�
��0���5�2��Ʊ��7���9�M��O�ĳf�/Aԁ%r
�X�wG�+,>J��6M<*�VMJuץ��#1/�*�_LQ��ZE�I\�@Fc���������;��G�@�� �X�m]�`�xg]���������7��"����ȼU�YTfhq= �w
�VV�o��:1�a,�n$�((5���TH�/uo���b;3rPCDO�W�LV҅�jot)��9�'q�ob`��������n��xH"��JB1��������WHv�#-�Y�~�0�"��]��1��H��:`u��_�/c�h�����u"X3&����ןf�+�Z������*���|�o��/��#�2� ��l����N��I)�g��큢�k�gՌ��&�Z�;�M�m�:�	�w,��d:GU�����/
^2r�)S�2.iZ�N@���A]�:	����Ş�t�켲���[S�rIDО1'N-�%�e�UIA���æC�X��M�ށ��f%>�	��
i�,��N����ӎ{y����rv1�H����v7�:�E�8b)�UC�/3`>r���A&(�3��k�s�=Cd���9g��D`Ԡ�{t����q�y�Q����L�C�w�L'�����M9����k:毥vlӤ<���*ZE V���tM���j+�?���}����EAA}��ũj������<�}�p�}�,�d�4 ���b xQcra��L�����^S��!��)�K���&� � >�8�l�s�X���j-FjF~���?z)�)���{���[�L�e�ߒ�!��������* ��H!�m����[V)�����?L�m�ež=B�<c�ㄥ���/�yFz-�=�TVv@v�3�������4U�r��s����tܮ����H�a�u��#��asjQ@EV��,~m8͌&=K(���zb�{]TX)b+ �P��YȾ�����4��LƬe��ѿ�]ծ�C}h_Y�?���D�h$�;&�2���^�{��p��}����w>/,�D�Sa��]}L���H���I�]�S�lu�~�����N�>�O�A0^�8�(0PR��g��s��A4����W�P��6[5��A��F4jr��	�7�dD#�u�}��`$l��E�AC�)�ՙh�`�n�/Eo�|��j�� �ANwLש�ct_9�<��*K�L�v�/Pn�i�~�1�^p��qy��OlR�ztu��RvnM_r����|)fE����o���p-_C�I�AC��H�hn%��N��L�ŁE35f~ɦs�q����%9?'�$4D�{`t�i=�[�i
{�k|�֘�M��Acc���.j��Q	�ȭ��^ E�3��q4����=�&�P��q�jv��Mߒ�����)���ʰ���7w#R�3�����N�� ��q�t*#��n�)� ���N�>�~��h�S���m�pHߕ&F��_�A�^򢽟o*�+��B�W;�u��a��*�uz-���<=�Nbų?"���j���'��W�a��\H��S\U+9�>=��E�qQ�{V�숕V��&|x�Ӭ�?�9�w5O
��(6{��N"�S��8`y�
�s�I��^�j>V-¹L�vx^�KFR���)� Ax�"�el/�ݥ��K�f�u��?����֞ZV��6�~]�3� ���ڍ���"'k��N��j������� 桡p�����J�[�s��cn_6f}Mj���+�M{� M)�'@�Σ�c�|+_s�4J�t#�1���O��7��%2���ä�/�����r�'��e����g��ժ&�8��)PW�qa%r����}<��sjc`.��ʂ���m3��*(�kz�i�<�<g<�+�F!ZL�C�+�Uɡ3��ᱳ�,���ܛRֿ���>A�c����ݲ�ϟ���bx���F[�ރ1�b��5�l���<e0�O��
��O;}c�LmI&�#Ѓ6�i�1���\�^`����j�2�W�r�b��uyP���=��O�KxT o��F,�֏�2�}����| ������t�4��XL\zS�QK�� 2i��%����y`$J���⮛���$	D�q�"��c��K����C9���������.�3��%�,H�1P;ۑPS6!�4���^�K��0<���^b��b�@�� ��I9L��R�L`X�yuJ��%Υ�C�� ��D�m������-����L�ފ���@Q��rČ��h�>�a<���b��c�K�-�t�N�+X���¼��!��3~�3L����I��O~)<�$��ؾU�|�Ȍw�2���GjT�	iV��V�I����E�H�`	�ߤ:P ����n'��P�nd���U�����T\C�[�v��|4q�o�Q���������\Y���G�%y'�P~��j{��Y�D^��W����8������R�+&���NR46i=�6�Z���'-s�A�i��q<�@u�~2�C("�W��|)=��YV
����<)��7r�3*��dn֛R���a׾��s/-��=D�W,~�w����2A�(}�Å�+c
g�c'��lR�Y�@����O&M���[�#�ז�H��c��b�;��_��@A��Q4oP&� �乄b2al��ùm��T�SՎ���h��&p�㕈O�5*|Ytc:�=�(cp�D�+��7`X�h�snj���D�N�,�Ί̸��3o��SB���ypD0�;�wY�rl���JM>��tN��	���z�a9`��}F���j�աFp��2N��@�3�F|I��i$K�?r�]\��Z����O3��_f�ךS�/�����rYu�|���|����wX�Bw��5��e�E��Q�5R�M^\�l���S=z���/�Oa�o���"��y	�FU��9����\��~/˘]~��1h��fID��LDS��W�I�uXp���-���پb���l#4w͈?\����k4ٱ>B�덿b�c����d 9~Em'0���&��[��ċA��=7�J�����+�~�/0�s8�ӣN�d��9�lu�X��{��]nv��A1���>v�����s�b�����ez()�% ��P�vQPb�����KIwb���ky�O�D��F4vd^A��#�9�z����=2]�*|�`��6�yT�N��|��ߨ�W�(�͹KYL���r�jg�H r���"l��*D�2Ml�5COAQ�Ӄ/�^����2̬#/�Ma�#4*k�4���
/��-�Ču�3!�R�1�K�X��n_}��^P�}�Bvś/�q��XӝJZ�Yik�G�����N2����J����īc\�G�ċ�.�K�C�́0��5���ᇫg�w���"�����ɧ>/oi	w����J��>��_tz�����ΡL�J��>^��k�I A��<�k�\��N��&�� ��M5�b���>]�A!�d��/�C��m�i���-W�#���Ak^��������2N�-�B˟�����������)�%�Bcc�<��}��wf��m�����@����1n�'�Y�k���T���f�>�ͧ�Q7��2M�Fr��|����n�0m���J�nx��z�N���ְᶂQh����襢zv�(}d�||����%�DZ�n�>�٥�F�;��������DH�|�1!S��y��j5@��S� �`(AȔ��m��'�D�������MW�H.�(v(4(��~ã<[��6��Q7��@v�y���2�ydQ���>��+��V;2T����~W��Nh�k{(�������J��H�oni�B:�G�^�ذ��
7rhy�����U��%��~����<�}�Wcv�9L��#p����6ey�?V%/w�۠����gҞ�٭�ݐ �N�n%ue�����Z�h�T��w@k���Lr���^�C K���K0��w����C�_��$�'≁b��7�Dͻ�97i�`�Q���갏l���)�������:F�u,@*�����4bg����&���k�����9]g�k�?u+4,(R������7&�,������x��}F�s�#3x��D?�/۶��<$Iʡ_V]ߋ�RIZ��&�%*Q�)} s� ?�Qs�I��(1��x?�[P��JI�?����SDv�_�K���}\4z.��������L��F���H������KWeH)�g��yPW��o~͠�Ñ����� d���C$�4�L���m�#�s]y�����nG#�FA��^�|�Pw�wJz%�h	鑭%+,��35���	�Q�Ⱥ���CQ���k�m����4��t�# ���B�Q�07
i�
��!�gfHl�YF��_d�9-�;���IQ�k�b��#�vV��tt]�'����,�����'=͍�Ͷ@�W���'� 5�%Gt���3p��΁�\��0�"�Sz ҈J?��~r��~Rz>N7��![K�կbX�h��W��ڋ���o��,:�y�A�S���|dI��ΐ{����t���T�����p�uT�-��F�'��0<2w�PUI�����ͺ	�=��1��P|=_0ʵ�d3�8Iz.�[#GŅ�ϭ�a�ڗ//JV����	T���I_�SX`���l*:1=�Zy�Sz�� �>�G7@��,��УAM}�.��U1?F�-;��:�t|B�Np#BU����8<�
��N)|�*�g�o�1fm��5��.Bv��	Qk~�~���4):s���[!��HI�� �/��f� �=�%ܠ�t@?`��:��=?��'�q.A��û������p��"Q
+��ͽ�uf�K��gT��N�.� ��X0z�Gl�
Y�z��� w$���#*}J��^���)�m�41F��{gUCQɥ��W�L�O�Od!_��H�=y�3R� ��S��b�8�� H}�7�%�>�UXJՓ��dBH���nǲ�S�Td�BE����|7D��c�{o�|�:> ���q:�S8G߈���"���2ik�Rh�7�>pm,B����Y��m�AQ�<��:FH`������Y���ͦ,�	�����9��r�f��$:P����}��nb��AL�3�o�B��!(b���&�`��WJ:Y⼉�#�P�'���{J�b�UF�)�}a��,�PK�낿uWc4��J阋��j�o�#������zjJt9����y3�F��t�$+ü5Z�d�IE(�. ��u������uǈ�:\!E
��W�$d�h���}�و1
X�x�]��d�����$�Y_���ֆ�I}��E|�ѾO��c͞�M�����O:�Z���A!y������߂�r�)��[Bղ��<���ֽޡz`����4|�w��Qndn�������m�X��AE���|���߫0PLY*x�*��M9��U!dī�x�;�عa�O~�J7�\�h�zF����� �/ ��N�a��ySO(�tN�60�G��q�{��dT�5���o�M�$����O
��5t���F�aփ��_�&�TC�������v��'}��� lhބ�g����d��5Ju$��,�} W�9���[#{TKj'��߮�$2�:��T]-߇޶R	��f�7*��%<uK�����,�e�,��4�v�)�Z	�A�����~|��fɩ��{�YW���tJtFm�m�˛���<7;Y����w��9�73���/�kb%�����y���c�{|�$|@��=#4ky�/��a���ʥ�Wl��:���-�PL�&(�47g����,~��GhP�SQ"�C6��7�cE%��W���}�{��|HẺ�s�Ȱ�Mv��r(t�tc ���HX���j{��=t����ƻ`�<����-�`�����濵�Q."�6T���&p�EuО���֐RF�V��M,
ߍf��"	�b�[Vq��²XIz�H٣-����0�_#�2�c��f ����jcjb����Uyl���>_Pw�y��8��ѫu#t7|SEn%���ߺyJ���y�M�ߺ��[3�@�	�bw9���*���yb��%IT����ͬ��T�@n���P��B�.�(��l���f�p�&)c�e���PȲ��(ȇPG�s��[��T�k:�?�N׋3���������׬ N�x��+��o�G��[������fAWOB��	�ҵ�\���6`���j�
F���k�ky�5p">���c�����Կ��oF��nL��ԟ����yeP'Ag�oPm�4>��bd���N�T�3J
�XϬ�N�-D�ůW 	7s����QDB<���x}c؛�\�E9Z���|��ŗ�-3I0ej,�L�]���o 8��"pޚ�#�!V�V��x_�5��m�ԠZas$n�4yY.�I�gs1��m|��?~���X�����?2����7�&JF�C�a'����;��͆#����J��)tj�����2W0݋g*c��C�����T��NaZگ���T�'�Jo��>�G�s<��_M�)���\��bMz|%���Ϝ�u����(�*���Q�J� g��e�w��墳 {���hp��j2ks��2�!�,�0wA�[���q;�n��R���	�m����I�D�ثy'��#ǆ���F4���x�UO�G���c��^�޹l�F�d�h��WD��Ű�:c���@�s_B`U*[�y'JfI߽��0b��h6�&��������5�y�����c
ӧ���e�~�~�we}���U��Pշu/�O9�iȌ%���c��(���瘫�g=
���G��7zL"i袲��qx
�� �%2���k١U._u�`D���_�'�|�d�XGM�-s�
� ��A�Z<a�tE"�l�_�F����_��9�ґM%���f�v;f�4��m�����B�5E� ���z�R����3A
5�6�?�"�3O�YzĽ����a�3gy1u�}�ͦ?IHT:Mz �.&f�*n~��G�F{|������e��Z�� ���ٴhu�"J�?�?86 @�,���]{� \W�`�kW���m�|:A-Amٗu�u��#L����#�}�q�$G���,��;_��7�{'Ն$!t���#�?��.�|�)�E�C7��J��ˎ�} �6RJх�Cv��T�`l��n���"";� " n�#�M+�Q�\�T���3���L�H��/���%�>��b_��wwV=�0����rw�L�GCo�z�[-SS*�*�|�����*/
$L�؂`���.���`�I�R��0���H������L9�g���bm\6,az��E��T����F�qh6�+��C�3�x`��/�/gţ�'�����8��`�}Z���xh��.��H~���t�΀� �цDM�X��]�;�,̬Z��K~�K֦�R�qR�W�,��;��
r&��ƒ oP\����-�,[����p��̀�V4�pZ���Ma���j�ՐhJ��r����P�F}�8�`>>����{� 0YD��o�QV�@!��ݓ�g�s�]�n�+鸈�X���U�G�3�f�6��)���W(!�׺�M_�1�?�B��w��mNX�|Mh����a�T,s��Е�A|�յ�iZ�[��Gfb�ɏ��}q����g�d�L�=��e]M��?�.ȇY�,�m�D�y��e�Ou��=�[�R9]�x]
��A�K悃��3�������*uC�>2����ۘmg�_]-��ڦ�48��ϥ������giP�(�'T��� a�cFi�D��J�R�C�!��7]�AQ��z�Qli�G����@j0���+�>1�&��AF����DQ��^�/;���&v���OB]4�n�}/�&�i	�+J=y��-��>��v� ��K�TNmǚ�x�	�}��+�*l��>#{��B�Q�*���N��|+�U0������H�eX�؅_����@�>�({^�8
�@�L�:��@}�t��f��7x�nM)���g���1�X���@� �x�ά	��p�d��i���U����k�?�r��S�*o��5L�JtC\��:7����oiR��lr� �x�ZY�E���r�
�yY�$�M��r��l�R��2jB,R�N�Zd��r�������Bg�^��	L�+�O,Y�̿�ъ~Uh�0�vnބ�g��Q\�YI�B�����Qgp_I��X�Z���Ǣ{0�y��OJ.���S BmQ��M#�7��^�8&;�LY���-�M�h�@�����Ԉ8��ί��8�6_Ǡ�L��<(�V�"?u	�Ѡr�\�diz��x���@���"AD㶉��䄤�~���Dý�_�	8����T���[@F���䖒.�c��K9�4u�Ex�nPߜ��D�.��K@
_LhU0�"�	~��R�W��Q��ܨ�����ME�'W��N�g`�-XJo4�0��0A��QD)J��r�)����NAo�bj�E�����a��g�)��,��'�?z ��Ͳ_ڕ��}P�f˂H߈aҼ*�V�"(�c�9�	'Dgg��Q�ϧ3n+M0��Q�}���9<lFZ�^��͹�}<H-i-�m��M,�m�����j��Ru���y�<���ϸ5�?��T�_��Y?b�p �Ik�e��_����(�<[��W�'�}f���9�L�O�KR�����h9[� ��C����G\g5��,���˄��V��'�!���;�_E65�J���N%�2�jˮ�	}13EN��/�*��۬9��C�+��A�>�n�|d�P�1�ӰN{!_����g!��y��bcx��^��S����1�^��BA�ψ�m�gU@`8ue�d��A*�5�"T�M���c�L^�@���@�c#,�Ŝ�Ǽ<tVkZ�?���$D>cSaf�qPn��~?�N��t�&a,�����8�zS%�,u�c�h+�����9U'�/��4�{`6��5N~@��7{q�����;|BN������nk|q����__�DN���KPED����ǎPˁz"Q��ߠ��N�k�:7��F1[�m�ҩ�uu\�� XRX��=�]!��C�Di�P�+�h�1�L��S!�p+�ၰ��������c�T'���$*P�i�v��e�y�j�7�-�o/$.ק��%��ˡ2I��f8��%� 
K�S�ޜ&��"^9��n�+�ȡ,!�����˄zf~2�5bQ�=�`���d�#����"��7��S�ac��å���5B�?��2��ߴ#����ZC�����_lS�qZ�[H���y�/��ؽ�#�;�4�T��g�Y���i��o?=��X���^��T�>Ľ���D^�'Ȩd�� �\�0:��٪	��$+��_��Xʍ���R���q��903�ERp��:�梪�zc�I��!
?<�>JTm@�D ����>;�����B,���e��5�r�~P6r�P��n�P2(�8Vjw����X���kǌ�Y�s�� c�K𸝷��l�w"���I��;��V��}����5r824��&E�;�ZN��8p�Ƕ\�|��+ό�S�a�I:��O|hs{����)�F��K���m�zA�YCޫs(a�J��o�s�G6[���
�~#�Q[�����*STaw����" ��?�����f�"���GR�!��V]|��e�D2����u� >�W��9��^̲8�1�������/�k��,�_B�f��j�'ĕN*���P�"o>N;�B�%��nfco+����bPrNo�˭��X����E����7�U�[�-�X��@�����/�d�XP���`�:aX���lj|�?�Ou�ӥ��4��a�.���[�U��2��u]愛3��	"+!%e��p���#� �D�y�G��Y�d�̩���+S��V��y���*?SM�a�K�1}���¢�{[��0��o	2�ͱ��WV�X����ap�!%7t�vjH�\�X�/yZ��a�9FO?�w:�}��+w�Cƨ���K�O�Jg�"�Y*��6|Y%)�Ib���o��^;�L��;��SB��K7P�X
m� �ej��QN�	4Uz�*����9����u
"�3%�4Aw����{�{m��*� fS�weW��&c�Y	x!�#,Bb�Ϊ�G��U�:;�����&ۈү5��N5>Τ�z�d��'ع	S;%d�(�,Od_��p�S�:׫�O��j�)�l�8��4ɻظ����@I��$>�؆)i3��Sո~�y��!9^D���lT]��W��^Ϣ�D�Jc�3�����S��){�����x���p�an�/�4Φ�Ħf!B�kW!��mO��-�ppݨ��k��o���JP��dvT^\*���f�زI֏�G<ՉзlGhW�8���D�-�箭	�X�\��95�+5����AY��r��Z��ZdA�s��.�ܢ2��
h�=
	�{�s�Ob�k����UΫ����y�`�ǣv����������	�W,�5맫m45�m��7�wP�Kl8f���V�I�h�3�G�b᳻I��w!.c~��/,����]6Gw�4r�;S������t��y�R���t�>p��}�M}���=.��Oo��C��J�CyͭVR�x�w��Hߪ��V_�c{Kw�+c1�R
�_mo��X9񿑖����EJR�p�D�;�nR8�Om~YJ��k�5�kJ���B-�����,H��N�0۴s����aH��߼J�T�oJ|��������|�����־�E&9�D.��?�L�~���p���]T�N��rw�E����zX�7j�Up�uR^�m�Z&�Ie5=�=��&
7�%s[�w7+~cԘg$�z���V�c��%�;&��ۉ�� �����Bm 	穈^��Fy>�9Bў�0e[�H�pC �K�ǆ�Am�;P�����Q�1����*�T��^����	�it����Bko�Y���?�t@_z[��=�	�D�/�'�?Z��~jI �צ3��@)�	fe�vm�c{�s�-��uz0�Ǻ��Qhl�1�=�{����o��Ey����C��X�v|"/�G���T�c���������P�2�rr�n;j�y����k�9��b.���5��n	8���o�S&Z$���B�R�RN_>�m7A�\6���Bz���w�����	>7��	f�Q��;��c�n�{��F��"/C��i&(*�i�)�%�)�)��jߍ��2�X����@rKRWJJW��Ma������3���g����3��|_��c^?��FGL�&�X�\��Xk��Q��@3�k0���VGE
DP=��t)������B�Ias�ӽ��ڍ��]
�EY�a({�U�M��8��?+�Y���x���&�EgQ����b��.��(���m������8Gs_�?��@���ԙ-�R�0C��n��iZ;�)�f� r��n�e�Z-���	�h]@U��M>ݍd���
.�-���x���UL��\��T1x�uqC���7�>WE�b(xGF��G3����rl������P�R��F�f����'bY���N�h>���ĵ��Xz���1m�Jn�[�q�tLL�3��:B�<cY� @�z�;o��!U��Yu!�;��i��O=2b�_R�؏N[��� *yuSZ�◳X'�)ړ��2q/Ca0q�4����|����fc�Kp%|ub�.$���PX<x������h��Z+Ԓ���>5��ب쫕������W��ާh�c/u�S���S(��5����ڛ���3�N{˓�L�Pd����yʍ�X�P���Biƴ�S�F$6dЦnk(��l<��t���'��� �*���]��.�:�#�t�� �Vϼ"*[PU�]=	;ݠ��Ƕ�K�����0ci�BU$4,�x�]"x_���zW��#�d��e	��Z�ü����ꡛwDo�0p:�q���m$��܊B�H�-�,�<�ޅ���n���yşBұF
��|�2�7�K:�B%i�d!�����Ӡ��G|�F�띌2/�(��0�¾߰��ӯŴ��mn]�:D����ɣ�;�@���G�`}I��a:�и���:/r��S�G��Zv�Y��iq����;ߛb���,���W��+��s��� ��!��ߵ���lV�<������w1/0UD=*�y�w��L+�����OK-ǁ�	�s�|����u�W�B���!J����Z{��`�S-�V�ф���w�SL2�/H��T���MK��
��;~�MS���JHO�Ocv ���T\��G��v`n���<��}����OQo�G��B����{a�b���F���.8�-;o�v����d�gc����:��U����t0��kTG> 	��E����6&�[��@o��Ϥ��Yv
����g��Gӑ�X� I����mj�"�5=���-��J�����K�����8�줾I	uȪ�gc����g��9��iа���j?�fۃ~��4!��^�̔g��Ρ��O�x�ܦK�"�^[�Qy�݃^��9�vE!��ח�fG�~Di�C����4�9�b�z��8���f�5C����hq���b��no�g. � �(��_�x�K�!��
By���B>�VM�eIS�0Z�>P�C/W�@%,<����"��D������^�8��a屩�����ڵ�LN�1�HE��ȕ�m���L��bX��W�qj�՚��"�ǲb���:��	�;��.��aOԙ��f�F�(L�����^�ڞ����.�cH��4W��MK�����j>*�&ۦ
�M�i<ю}���j�
)��1	|>��~���.W6?��b_[Ǫ��z��ұ��
�Z�n�ݾ+Sm�����HXS��QT[kY�	�YC<���)���{\��薌�T�	P�p���B
������H:JJ����r"�7V4z�s`��"GD�Js`�5�1�ңq�A�\[�p<�h%�,JD��6��.	<�B�i۩��ͥF�ɡ���	�]Dz�5f�L��C?�.0M��ͩW���-{�0�r\ ��,ғ�M�$���{�;�����zW���j�;�)��W��U�����������3�d?�i{���;�auM͚�Q�TG��+y�� &U
�h�+��$t���̶��GǱ�w�f�4��p���l��;p]q�F-�;Ѕ�78�B��	�� �˱˥�_j��wC����ߦ���^�9=�'�-/�>/Ɗ(C[���7���tt��d?"��1��r��������j���ܗ%�b��P��N�<���4%�S����6�� ��M�_���>�6��?���f�`G�[��1R��,�`�3���I�)^p�F=~=*К)=��lz�`��M�&X�D�beJ,�y܄��Y�|V|��f�hn��ʣ�n�����(Ι� ��	����L� !
��iB�U]J\�=����c	,'vF���x/��'GrG�b�K&O_5s��+1H�j�WL�bX��6�f�5N����Ĉa�C�g$ɤ�v���
�[]�#e���0ss�pD��p�GKR&q.GL�V&*��1���|B�*N%M�kس	j,̔S�a$��n��Z��z���:�N�uc���|�I�݁�t��@�^�̀+�0����i��& N4��+��qk֭n���F��QH�k2�y�����5oc�ff�a^)�,���
�d�]BoE����é/����J����Q�f����
	�b;��x��J�Ք.��Oj����ع��8��`��n��N&h��$�$�ׄɼ�+K�#}g�z.�\�D�&�֎��sPi�]��>����U�[�Z��4ҏ�"!DƓ0�I���f�1���ʠV�V�5t,
(a�c�E�ݶ�(`e��o�g��L��j��ɛ´�hg�"&������Z]��&����-"��Gu�QnW\xA�Q%r.�s�^L@EG�ҵ�t/��Hp�R���Tb��T9˰(�����2����y߫�����/���j����'S�3Z�/�1��C�-�ֶ�:�::]{������'2B���^&�V����g��
�}����:U����2��D��΅R�����4�b��1��Xc�6F�w��U��}��P��}Ԭ�����IJ�:�~���MQ�C]��u�|���f�]s���%�y�_h��)�R����e�rO�G�Pmm�ܘ�H�C��U�����i�?7��-�ȵ� 7%�O*�KN�P�tV߻��"��v�*O$8���i�v'+i�����U�%i3࿓�G/2�����ĩ�Pv��D����,"�k)+�y��j��PK���O���Y�8?#jz��	��G�Lfe�w)�u�~�f�F��"}���^?b� ���ߍJ��OTeι�j�dI���e�9j��28By�8��ߜt=��kSX���/�J;���1����2�S�
,!��÷�Gi�����L�=R'W�@S�JJ���*�o��6/��#�Kvr���UB�����?�$�AO~ko��S��WݱZ-Q��{<�J�mjrt ��űM'_e����yt�Z�눅&d̒d�f�z�4�%��fܛ��n��fu���bG�")� �k���0yK\���`�����~�$ɘ��-L"��p��n�;=
&*^��5uw��&�2\�@�k��S�t'��ힷ_d���a�;E����6h�6�_E ���Y>�$�>(�V��[����7u����
����9��&-�����vI�s�"�c��,�ݞ��2�8��`���9�:I��	Շ� �	�t�4c��I�"2(��$kqu#F6��F��(�M�0���yE�� �S�P�8V=�T�w ���.XW9�*][dI���@1��w��U����b����p9�˻Tv�{��n�I��[>�m��	��i������捥����7�~��<��Q�S��HJ�PF3{v=Z��9̚��؝�&�Ӊ��o��P����B��k8Vn�V�b��֍��k��僈���6MJ��;���8��*f��tR�y�q��������I�S�]�Hmkw�蛮jwq�!e ��;�)��n�֜N|�׸���G���Vu�e-)V�|/�y����N�)]@�1��C�'l��=�҅b;�G�c��>d0^~j��pd�/�p6G꘶�1�ō��I6���Z��q���WuM�,/ �J?v�e�����uڨBD>1 ��ݜ�?��3ep��D;w����)�B��n�k�5�G���#~���b����ƽ+�����R#a�F<W�y��7e�nɄ�`�<�O���MO���P�N��B_�`�c��S�#%,�K?٢fWhgy�v�]�����,�@<��;�ץ�[��Ϯ?l��g�i�+�a��A:=e`�l�/:�ޓ���}Uj�`<o��uK�+N�sr��`E$X�abO!/���L�o2���2캆Wr NH���M��7���K=��Yc�%f��Z�ܴ�>��@zMM|Vm}E������ա�F�L�(�I�Љ��L����zt�b����y5�l�e �W��1b"2�^4�G�{��P����^����9��A{��6~�w|Y]R�B��O����6b���,�b9/3��w�_���zJ����+������t�y�JǡH`bn�2���T1
}4��H9h�Z�q��VpD�1���q��0�k�vQ QŅO��������#D+�b���Q4��q<J2!��ܵ�J��l@����V�<���X�T���e��;�)�oɷ��[�cѪ���H�x��]^B�2Dog`�p�Jz"��c��EC�v�N���4�X�%i����z�P�����1�0���CB�Xq����88�ᕌ�?����Q��8�s��+��] ��/���9���/ �z���y=+�Ntא�$$VՒ�=�:%(t"�cXM�c{�$/'a�dY
���fГV���s>��ڿ�|{�	�����CM9�W��*��$�&l��c�Vp�(o��r�T�)+��M4w�/G௧�,Bw0���~]Ey؉�0~��^ ��)���b��k]�Z�U9��)�E�Edl��
����w���Ү�k��y�w�xd�%�rCk �����F�`��wΏ3},6�ϙ���2�(|��l�Je%\��z���+��\"��m�G��rq��I��16
����h��Da),���9Š�<R�R���n��\�Q�S�8�qԡ`��������aJ)0��aL����.�C���/$~�m�ZC�d��p�IBh�^����Ph;uy��7���r��7b�R`/�3Ŧ�`I����
�;��MT�X�.���͞����T�giuɡy<0s�,�p��3���s����׉�lK�N���L��*.9)��PNT���wZ��!	Bn�͞r�D���"�(q��@e]5��W��Z�_+����i���!���P��$+Gp�\*����ܕS|I_�S�(n	���Y���`wǒx��6�!�!�I��B��-q�by#���u~��4M��u]��?_j�Ɔ!K6J�+���:�Os�Qrx
��/�����Zo~�B�J�a�s��>���XT8���@�}��O�=*�$JAa�����5'��z���������[Yӡ���[$�5;{o�,�Z��kU�S��G@�����[�`����զ�8��1a�9nJ��l{;��kjkTx)[�ǋ����Ϻ>T�`[��C�ݥ���L����?����?]����A��9M�3\Z�%9"���κ/ в�M��x��u5���:��������f��ٛLz"�h"�%k~,�D��+���f �U�z3?u���1��?B���rR8��|A*-�;�VL�K8�����f������:,j����e�I�Sq�u\��(T���Sf��� � Z�y��J�v��,�K`4�E�ÿ��I�Q���	��㗩�����}�0IE:�B�2}f`Nv���:0\Ѿ]/V��Hi���h��
��4��?�>s�GK����A���:4�u}B6|����~��)���n�E�G#rV�F�%c}ę��8���83��j���!���TV¼�6C�cL����6�F"�5_�jP�̓Uԇ��ٲ+������-Z�����I �\]�N0�m�J��_~\�7z����k�V�}�؂��ά�!7}�f��)Y��7~ډ�"�.4[�bn��E�=`��Y���s��^�K ʂ+�_P>�^oZ�a'C֝sΤ
�i�r_3�W6ə��d;�0�=%g��B�tp"[4q�D ��.����꒽��@;z��r�l�2�^p����O:�Gns��W�"(�]���K���L��(�N2�DC��R��r�*�r ��kɬs��+B��V��w�����m�!e�����bd�7����ң��f��_"�ډ"�����k��Ah�B�߭B���b7#J9��F�o��T>F�A�0�t������esRDr���<k�A�`g�{���RY�R{V-yT�#���c~�u��V	��j��M��^V�&��-��>�uy�vF�D@�a_ƀ����Gʚ̴="�f�H��'�k��R�l-�?)�/�MoAK�{-=��;�!Č���!������.���r����(}�w	���J9\ݮG����(���г/�g`:��J.V�, /h���s�M�!J�G�S��N�!��+�>���a�e���S�3��Ղ����btlq0,8��/�Ͱy����)CP"�=���+�Q�<��1�@��+.w�*�-Ɖ��	���mB��b2�5iYA�l��z��(hf��_�=qL�;c�wE)Ǫ�����k��&%q��`�U�-�	�4�7}7�6�m�S��½0� _q�O��ϴ+��!ôÿ2�~!hC�S�RVG*�z	�أ��,�}S_��X@�����A��&^�G�;m�v%���Oä
��º��u�:L)9�� �B�p0��r�k��EHq�����&����p�=��"莈����u��KS)���0�7 �6L�a4W9�\�Dd�������}�%l�6��!�,�X�_��xf�Do��T�W�#�Ne�ȷW5��y����e�?7)���Z�>.����qif@��R�S�[HxF���n�E�0]�u�%i���pi?�H�u?0	��_�oF+�:�w�JfW�����qx��އ��%�>��� ���z@�xҜh &w;>z��Zf�����/u�Є"�����I���T�-Y!��z�{��|��c��*��1�Z�p��~+O�`��0��f�E���*����䔣'�z��l-�rB��hQ2R�|$����-�J�~`|�� (O�����b�Z�o��|c�敱�MA�������'�	Kw*��-���@-;19�8����6띊��TSz۹܁8���Z�%%�h6a8h��[�T��!2$Q�4 ���s�"���\�B���PLȝ?u"�vJ�×�T]�&��J4�qٓb49�>�����;���Lnu�(\�uܴ�ndg���"1����Գ�x�������&a���zP^��4E�~H~��kە���nX�f!иn��ѻ�������`�����W�ߜ�8ς��*e��m�.żӒ��d�Q�Q���]#ݗ�]�j�K��%�PJ]�KGʣ�-����%)��F��������0�jp#�\���u���[5���*2o���w��[c@���#�[s����aӏSe��<]�`D��J��_��8#AQ~�R���4�i��;x�Q�^YА� �p�13���&ڌ�-��3}NKO��f��C������W")�,��~�� -�\
驼��Un"z���\\��^�K���}8&��§s|w�"慱{[���i!�0Qr�32����a!δ�w����(�5+_�ҳS�.�H���*��s1���!	�9<��cw���d%���k��	�\J����#�K��1�W��Pb���{�'����ʱRj֢j���i�o�ι3HJS����+��ݍf����gJ����e��w��q�b�ʒ��jPa�!G������c씥�i��0A:�(nR�8��Y��l<��)UT���WO��%�%��+��hg>��G���r�OQoͶX�}�ҡ�^]ٸ�~���N�Y�C�G頂�s`$˲O�3?#��hhk�nJ�WV�GSF-��>��9���~j��.���u��F�j�~�<ضM�S�sF{+�G�����?��q��^���*W���\S��6,��hW�܄?��`˻s��E|6�{��� �_}��2ˁ�[(���٘-��ɍ_2)�Kʨk�������R��-��j��Y��-U�H���$� <����=��ٖTjG�Q!�;�+C��jц�&B7=x��dz�4�3;��G1�������Gi�VD�hL����"3xxR�1�cԤ���ʲ˾T2���c,�������IeO�Q��ߙ��&��Z�X�3�����!��l}�/���z���q*�Jb	^|�����p��R`��8k�p0���'k�!�w�oc�,��FF%����vz���(�>�N��$���nм<�b��0�wr9)�ek��׃+%�ϵ��s���B�:���1w�U¨&�4�}N2��;�~���Ve�sO��˯cqY;�u]���L����9���=�kۚƦo2@�9B'=\a���v#Q}q��u]?����3��M�ֵ��C�K�D������^��� `	qu΂�U�M%��p� cs��R��f7�**+��l�Ë���[ݬ�I�[d����LJh�������j�'��GD+��{�R3 ��zzU�ĄDi:��B��:9�~�B�f�d�x'b�O�y�^C�_܎ne9*����;��l�Vp�P �1Н`G� +��Xj���+)��4J�(�s`�o w(GN��݌�������M��`E���l�+�̇��n�[�	r?��6{:�
��uⴖ82�:���K47�>�ad�o��ˀ��W���~�Z�-Mo��ދ`�Ў<c����,��Q8�{�._�e)�bA�	�w�B@�E�bI��[���.Y�-�/���wtW�D��u�n��\	���� �<ǿ����$�+��و���'�6�#��.�B8�X���BK�8���hz�*gA03����]��c�z�FW�&ѯ~{�V�`��;��X�;�H�!��:�yD�MjB��U�ꖷf�&���.�q��C?��]x��F�j*N>�wO�v"N@d`�ߥ����O+��Ǵ�uN�?xq���������"
2Kэ#u��
����=h��֮�VS2�;����9
���ݶ�.���Zl?�Y�7 'V�n�v�}G��<���³�R-��/r��jS���s"���h�� �*�]���.�z�:��������,���O�1��Yj���Y�Û~�q��G�)&��F�8,��c/��Y�z��kXt���whe�ѭZ���t����{��$�\�(��J�Wt4��Sn&��1��5����*^�`��t�7'�
���E)UN�z�os�X'a�o�)���6�1��N�;�h����D�j�C���Zjң!�&L��t`E�nQ������w+Yk����.
���	�R�W���*��õ��H|1>}������q��	8�4 HrznH�O:�C�Z�U�����\Y�, wV^�[Jנ�Iֈ'�GЛ�y��d�,Z�a�yLɲg��ڂ�����8$z�W/,�5I2�,�|A߬�L���٨b�vOT��	�Za�s��n���11Ƿ�C����.ޭR!�:�?�e{��4�8�S����E	l.o�S�g8���LTҨw.��}�*A��q�{pL��O�mY=WА]V$�\Qp�qb.y#�V�S�@�Yn?(COv�a�*�^{�'��+U���q��Q��qx�Ϙ��R	@>8wD�狐IB�dl�O`��C������n����k�F���W��y$�f����D��I:/ X�6�7�kZ�{��xƑ�0pr�|�H<����*J�9Xl�lC������6C�#�t��KT-�6��`�eY�F#έd�o�є�����PsD\�7u�hPnı��o�ճ����v³�"<yX�Z�ֵ<ۂ^�N�J���K�F'���9��?f��,�p���C�?p�Ia�/T���"8xE�'�^�K�mhs��(w8������L���t��
�IN�߄�"��?�R�)�5��>�^���[�˦ �e3����xL��n��w��l�6HH�ݤ!]+���:J�eX2,!�z�tLNa�a|y&��49>r�L�'O�h�7Ҟ�=�V Sԕ��޹��3�ӂ�5��ӈ�	���*�8r*{{Đ��X��o˭�����(����w�5@��a`�r �r��&=�J4r��M��iꖔj#|R9�{�Kwf�ww���Ԯ-���c-݇��f�8���q���Zk
�$i#˴�[�.���!�Y@��m�9�#�[H�`'"�qUCdT{e������]���m5\cy�D�_�������*���3Y�^d��T��
_F���o:�J����+o'}�"����>�	���9��m�Ðf��0�"��~/�o+��|Ad1��*�Y)vl�ꭿ��`x��,�)�$/i�]Y����Ǭ�y�(�O	k�Ǵq:�i���ڼp��o���������/�Rm�8���(���K���H^��>�1�P�?f�
�n��p�` �FH�V�����	��7$��w\���VFz�Ɗ�`����	�-j����k�(혩�K%�H]���fn�\�Ub�}r�do�c^i� r�.=��� +3�z�zd�LD߼��S��(Zkm�펩k���I4{�-ϐ���npcv�kVBn�褚5F�:�1q�nZ�b�[
h�#�z<��/�h_}�ǲF��x�<P���Q<��/72��M%�)�J��lZ�2p*�Fb��ͤ���Ϗ������,��!��K�i*ǃh%����ú��Ɏ�K_�9Y1 ���s�<1~8���`�z�z �f+W��L(�vk�7�dj۶���1d��D�M��eu\��ߴ������rҲ��i]���Tݒ�⹨�p��b#iq��?�����ۍ42Gx>\���Zc痸�q�B����.[��Ӌ�Rk��Ⅹ�;�{k)7�r��D�`���6�+�(bm���5����W QE]0�L�*h�^�R|���ғ����P���WG��޾|�)X�k�E�c�44��5 @�xb�8�J��ɕ��G�Sd{����C���ǜ{�F�k���3s�]���H_-���
��� �[b�;�amY�	>�k-��Kkr#36c�ҧT7�_�_����!���py��9�]��m��!�"h��|�|�{9�����n ��j�w�Vyl��9X
����{:����EG��D�Q�q�a�It�'A�
a$	s���wϕ��pzEE|<d��oO$��j�	1�뀬�
�~���K����b%:��My5X�� ?Tۜ�x���겞v�r�L�D^�5c߆��7]���pX��xv_�a�I�������T����;r5܆��a�a�?޿`�jYzr�YG����*VԶ��)�������x���WD����ܜssy+f����8��SwhB��.�'��Q�w�|�K����8Y�ɡ:�f�eǼx@P:��g��F*+�=�t�[]�� ��r���x
�6n���VhT��F�	+g����d�'_��/����7$#���fǣ�K �a"�������ȕ��^�H)f���������W��O���E�7S���󿤉����SJ���zB �d�kf���&`y2V�ǋ����&�~�r��9�<� E\�{M{��!��`C�� [jK��֫h'�D�MB���`�H��FM�^���x�-��[�����o!�iЛdX}/D.'_�`��E��|��A�m�t����I8Xv��X)���Ј�H쑃�i��替˖	._bD%>�Ъ+�ӡ�UC�_l ���KU�69�IB[_f~�O�����^��Q� �^	 ��pz���:�R��%#O����+��%��A���ļθ:����Hm�짼Su_���$����ތ���y�A������
�JIQ�(-�؊v5��W�S\H.Y�6O�L�� �`��޾@�9����͵Æ�s�|�{!���,�Zoѳ�r��]���[�ko,^{i�%�s�����Y�LR����K�m\y�0��v�=[��5
ќw�h���
�%���+���^�����/�e�/Nӧ���}շlڲ/e��b;=S��.��`$d���_-l(��(=U������?ޫ]+,��u�=8�/�7jCO⾉����X��$6��X�UGؙ"$�,|h}�wϹ%�{[ X5��æn�I��߫��)9g����1v�n�)��H�4�OqȦ��&Sʥ�Zbn�5N#�Cm����;�k?�������Xƣ@,Q]f��mhrb`x�Þz��#�@pr(�qlq@��RV�C��{�-H���*%`q����4���[�h�{�ŀ��
�q������/M�q��S�q�z�~�b�֞р���8�����TQ9k�E�i��a��T_��MC���j����Ӳt��#/h�y�ן�������u{�Ꮙ���ڤ���|��!����3²����tC���G�Rfzx�M*c���<�+�L�rb3�z��S�bo=ׁΥeh�(7?��+?x��&�&8f`'Ỷ�r��D�	�~�j��z9��4C��������~����_c�Q�{a�-��Ό/��C���:�m�F��ӕ��R��޷0}�?�n�����@t�r���D.�#�_�op�ך΋���l�_��x�q�Θ<i�4+9N��X'>q��Qv�~C���]�?}*�'��b�V33B�*m���l�6bL���i�C��o	W���D^���|:γe�UO����7!��R9G����Yu�P1r��*�m���^P����H�����>Aת��� /��W3��ɏFư��F��~HV�_C�E�J��/���5���9�Zu�Ik�lQo@Ś�ۯ�)ǌ$%v_sZ��ϫ8JI�B�
���e����~��u 2����OZ���B���vm�`p0��(=��,P�����%w�n� ��E���1��Z�����=K<��P]�?C��"�``�&@��k���T���~y�4�s׮Lʣz�`W��~fQ:-i�~����pb�>܂��LeA:���1M���+�N-{ĥ�ѝ4Kw_�/�[ �.�g�Ő����'ސ�OC�OL��
� �Wⳕ_Ҽ�5�� �:��:?2>Y�������挛�`u���Xg��.y�2���̖���#��D��"���4K7>��I�o�C�⪙CB��Yn�H�� X0��"([��̈=���+�d�ﵷ���a�	�{��ohM�`Z����$�!��U�c�F\������݀t�X�:J�&��� r���]�D
��~s�ؑ��O5C�t�j�39s�҄�ɸ֙��%}sN��N�/,�+��w��ڑ�Sj ^��l���(�Ŧ<j���/��l���GoVFk��;iVki�Y$ �0Ƚn��G$߯��A�ɕ�9��/�O����W [nq����c.���h�?nT�[�ɷ�������Æ]���"0��lj2��&��Q$�d<A����S�w�9�S� ���ǺnݩE&ƿ_�¯A�A�zH�+�҄W�t��a+�ΌǛ_��5�ژp��nW�z����tM��2D���l��X��F)VO���m�9���'�������F (;�0��1�'5T����e�T+\6�I���v	�RObDM9����y&��������v���_o�<bR� ����P�����Z	.����=�O��:�褡oħ��΃���d��P)�U.�K��t&,�D�:߲(�;�Ǎ�����'Ħ��*d����lh��x@D�1蠙3A?�D���]���.���7_#�����זX��Ps�UC��!5��Ae@�6��
���"
�m�c���ɂ������JΠ3t�L`�" WC�d�5��0mN��&A�J�_��2�L��+5��	�\��^ejLh��i
Y�(�!�������56pjNX����a�0�7���s����I��Wb�=����7���P�(��m-h,\�e{Y�}ҹ�����-�$m�1T�@��O�i�QdN�)���F��ɍ���=b�7
䡾���d��Z�9�"���}��+���[q��!����c'��i��/
nsgh�B��{V��
%
),��(~n�D3��+�_d*rg�9��3�|�.��^!)i��D� C�/ߠd�D����G��©%�F�s���u��;�e/� �b�E�mN���'A���ゎ^Ob�l�ΐl��=�~�i��!w�Ӱ{� �Uς0Cҿ�#a�f��Q_+�^b���"��p������d~�ynu�r����jxd������R+��\k����Wީl�߽������
=�Un�.o̤shԾ̥��O�XLv�q�q�K��Z���E�i]�B�ƃ�3�]�&��۫{0�{t��SÐ���&Dl�L>�.5�|/!9�8���_�h�=_��jP�k+<Ie�.5UdD=�X��<�9c9�ή����l�S�ӏ?����C\�S�i�GL�XVs锛6"L ���{[M72��yXD>�H�����S\�	Ğj��z����/����A���ؖ�f��7k`�d]yj2�I���!�l����7��)
��S\.�m����6sE�sh<0�3��M�r�#xV�E�P��dN>��&��춌���۰5��|�d)�53{�Dyj�7���j��$*�D1�+�+h����&Kx)��jK/���=���|"݈2�[^�{U?�;�o�0���4We���ރ�Բ�ͯ~���� �(���N��{�9O�Aq7�I�8/�_���e�II��,�]�$޹�'pH�z�k�q�?K<BMi?�\�p�P�X�ݮ{>:Q�W���L�-
jd+��s��Տ �Q����g����y"c0�|�̛K�1Ev���)�%&��f�4�jPv�5���#H~@�����8�XV�5U*�������4��5	%�?<8n�P����T1�V���,�A5Ԥ�����#<��B��;Lʪ|��~	�|���Q���B�Y��)�Z��#��B)�!�Y���q�����^,vC�QK��1;7@�O�	��*�E�}��86�O���`������Ǚ�n'G�o�F8�/�� ��KFu]h��Es�-#�\��s+v�h�����߱���,�n�J-�ӵ�r�����Ri޷��ʐ�0�Y�Hh\{A?[/K#҆!�y��)'Ԛ��ӊ��}.��Ձ�s�2��g� �� ��y�[yd��:����Q;�"g���1[q�Œ�U��o�(������;�&QNX���F�ou~x������r�P�hrm� 4���y�~���|��U#޲0��|c�fÀ��5��S��09.ơR(x��^6�E}k�d�U�Vd8�o����--8��סG�����<��4mL����%y¡�X"C�A����`G鯰3%�����`����n��~�5^4�����̑�s�6hE�i�m�7�[����J[V5D4u��߬����-�¸34@L�B��{���ɉAU���]_�Щ��Q�" ������Q4??�8�'�w�"S�L� ߟ�u��җv+�a���3��ļَ�LXmf����!�jib��RLCS��۞�S��}�F����)��� %�NR��A+�%�j���)���ZJ�P�L/�Ŀ��|=v���P�c4���� �il��d�S���H�O���v����2k?��X�|���U�Zu���I=HR"�C�Q�YY��4l�lN����]�y��0�v%ek����N�EI��q��3���5xmق.Z�6i�B�~@��G�Ђ0＀n��)��)�����k`F�ƚ�g�d|E��ed�_L��?>be�q�Ju-���V�u "]��5����QP��S7���*;叹�xo�s'�jgАe�s�Gu]��Ǽ��d&W,YIlv���k���Lts�{�;�^0m��w��P6�a.�|��{I3n.n��3�O`���R]:�A⾝"���Ms\_���r(*Օg�s�'������Ơ�1�� �T9e�Kܪ�Z������&���M|Y����Mh޶�O�L�Ͱ(,��3`j�����h]}9'+�ԙ�.�� �W��D��vc��$�16d�w�{��;fn��9�޺����������ک��	���Y%9�3����gD�K؍�>F�D��Þ���f{��^�'!! �,�!$�)ZR�7-`я� {X��g��A9/�]��1�!��,� ;�'�/�w��إ�̜f��A�r9gj��7�ڳe���c�:k��Wi�ќiI�M���%޽A���C'N�b��O�d�c?F��r�ɢO�"Sڴo�x���?u����g��c}�d�|=��p�U�*\�_�>��H�O�S�xOd�El{��uw)E[�z��գ��#���KRv�m2��7-f���'����u-�a:$6�qP�8��o,/nb�֍%T��{���T��i��Ѱ�7�4���l!���x�w�^T��5$F�&Zfc��kq��b2.�.h��+r��sfFf��ɿâ}�7�L�!�gڢ�:)�ĚC/�R�]j?�Œ03A,s���>OͽN��ᷝ��/�*\�#B�f��i18�R��v _.�}R�!!BZ�5_����~3Q#>X�՜���oR�1���<��x� }6��̕���It����f��/����4�����<|g����\ؙ�aE9�9��V{�X��#�1+z>����dՑuU+@0 `#�.�\8�ȷZj
Eš�R���f2�Ʈm�\�FO��b���mGާ�e�X���!Xava �m�:�;i��!c��o*g��B�DpH#�R���*o����H�������7*?w���*Yx��R��qarg2i;��0�~XG�N����>��z��j�%��="��ԠTe(�.t@&آ�ߤSܤ����9�=On�ݢ;���x���#Y�H ��o�	K�G�E�r����ӗ;Dd��D�3�u��p9�W��?���rcx���֨Ώ}5%kTMq8�Jd8_ς����� ��­)�-_���T;��۟�cd��Q	�@A����?R��M<R�X����CW�:.P��1��z��ݪ����mF/�u��`B�r��P�,|��@'o=������H��r7����l��Kl���7%c^��י�TWY2��Ml��{�N�|�Tx�+�q|���QN�:�z3_��e�(�3al�&x��W��`R�ghE]�z=��8����!X7��
�iwB�J���C�<�;�W,�ʒ<���}�<IA��ESk%?�VLW[$��˰��>f�W
fN����[Q��-?����FA�-�O����я2�B �(N��<�:ʛua�?{�
XS��;֡g�D�&_�7�\�9�*9����9�"�GL�P��h��� &�=��|�R<�[�=#��6�<��
��*���oP�WAZ-���h\-����1��{'"r�+lӿ�"��#�3;�� ���� f�8�5zM���5pyT)��̅���3�]`�I^�|�:�h�1#H���-��;�'
Ō�y_�yȝɌy�ѐ^,ii˧���G �Cھg����*��H���C����DmT6뛒���H���O��Uu��æǉz�P�l�ZS��W[r��+P�4B���@l⭃�_� G��4?�t��wS)!e���j >c��f��~����^찁H��{&������X�^������C媘���P�i�� �#�f��!ns��f`]2��5۱��ccEc�5�i� ?e�+6�ъP]V�
�S��@]��u�5i%���q�vP�C��ZM��0$�ʪ�N�YPe�q	���\Dx���t��A]���˚q� �N;�Q�6b�b�+8Ƃ��xn��Y'҆�5ag��&|n�4�Q�~�����������W��~���M��+�_�n�Y�tg&��T�%�Q���mc^D,��N�%CSJnG��	���K?� ��Y����Cա�}Uz���0���E;�fGw{~N�ޓ�,݉o��4����l��j����o>EV���8O�ޣ!��iA�-�B�;�&h���kx�7�&{��&.M��e�n�F��xɅyq��������W��|�K"���_}�kԊ	|:�O<]��J���:qC��-WN�T��AŻL�i�)Xt���� I�VCM��u��1o%`2X�p.���3*�ivZEw���<�Z7�:n��}�/��^L�8P{A���>Y�$r� �9!~�y���Z����;�NX�r;�I�U!��K	m$d����Z�&�!�uq��k؜&����x��;��{4oV�쒖6�2���u��;��u�ؖ�?^�_{��%׼��iUt�f��,���F�֨�P��Eq`L����ݤ~�}WE��7�����n�]�O@8tG#M�����=q)*V*��R��u�;z$��pW�+W�r��!M�t�P�������\��C��1��m���z7�(�új��O��!<����'������\=��5&��`=��%���E�r/+,��O���i�����%}�nŊɁ���ʮ����2��`�2F����O�NMy~E�ͯ��dj�޾�%����6��j9����5~;Qs�`�+J�c���Y.��H{� IJZ|� ���s(��P��OTB�tg�w�ȷ0��Bd2{ˑ��"�~��00��v�:�����^[�J�K�����oщqLP<�f&��" ]���ɂ�Z�����.�!��{Y>;��� 0xǸ�&�L�/Ȉ2�T8���K� ���p15jQ��Y� /w�<�`v�7����	dP��
˿��02w��9w��͟S���NS����gLN#�T�~���p?�=D���:����=4�l- GH}rr�Ű RVh��3	�r�Z�yjԥ�f=0i���.�Cqrc鶧�u��%n�W��
����4�3a�F�#���!�m�'���P�x�ުy(����S�V-�O��߮�J�oUD�PS��T�sY��"#�J�R��� ��y;���������7b1��@EG�Xܛ1�جop�g����y�������d+RE���Q�z���	W�mQ	�´�L'~���
l}��ٔR���K39�`��ɏ�l�78P���b��*z6���`:���?0iΌڷ��(������쁱.�3jb�\���ʢA�,-{��N��0��W�4�A�ŋ��L"����	q�/����
/�>�Xi�&F��8��v:��(�%�m"ؤN)l�\�$�r�yi�҃�p�z��H3C��`9��q��s�F��3v��k�p#z�yYǙ��Q1.�Y_̡��p+"�+��f��B��r
gW�᫆�d��ضi�r�a�c5��x�i;lʏo�-D*���L}Y����1�h�@@H]NZ�pAt�!�?2�)������q�ë����e�obH��,����N�����Ł"�3?T�4D�I�4Qa��b��7S�f� �\���#%�^�ʅ�	��y�4}r��.�ܲ��!�k�A��ހ�5�Co� �f�y���������)r�����{�Ѵ�]2� nD�9�/�	��L��n��\��a���Y�o�iB��t�S�y�.!������؞J!�C��_0O���)sR��xx��q8���<Mo���^rT')/���]!��{;fI��02(Rq)[�I���_(�H	pIsI֕�rۓ�ϵit&l�p�ⱇ9�#�,�1���_�;��V�|.v4�C��.չH����K��*��SH��9�a�h@��4�.�i������'�V'�˺�#��yD��֥K�
W���('�<� �� ��kǂ@�u�z��e�Ub4��g�cƁ�Q/ap:D�Y�pR���6�� u����;:�V��g_�B��Ɣz��3�:������P2��_DDs/�Z&�X��q���2*¯�D�E��dث &(��QF�E��3���x��V�
�Wc:�����V����Ѵ^B]�t�C7��Gai>A�����m%�e��@үI�\ee�7���b1����:$g�RA��aۥ��s<���#�0:)ӡX87~�k1*"�<��,��.�]���	t��$���~��ﳧJ����()N33�-B�33���lA6�&��&��.�)w�����I��p�1�D�m5S�;7L�����	�KX�ڱ]-;=_�,�d�A2?�������o���)dN���t� 'z����Aa�E>혫���9�}��v������:�/�%����q���lP�:Y���\�U�z{��3�6B���==��d�����
��%8/�]����&2Yy5�Ժ���rn��!]~GI�1s�R�=<X��'���jf�4���A���d�
n� �i��Z!:T�?����jl-���I�gK=���s%�nߵ7d�G2ݘ��]5�Z��c1�XA�F';���͠�Pk���0�(~�ǟ�El����~A�+R��P�l�����)�;>| ft�Mpo�H/9K!���4��5����A�|�i��[Q
��A~�ɝ���]�R��S��lQ6خ}���+Yv�qS�]�cD��o�,��X�:��J-�s^����- -�-�J��Š�`�9t<���mS
�,SR,��~	��R�W7����G�G�N�r�f3���%��_��4uqC�gևLS���}�����g������+��w���ȡ��>.�m*x�=+���K��������~F��Wd�Ƞ
�&��!4�T[��!�*l�_��\�w��j��o��A�$�ѥW���ڎ��#��� ��C�M�iAL.�G���x����U�hIh��(�)����`�����Ze0T��!�Z���u��|f�(H�!�EF���<�@{o !�%����BE�W���1۔Uט]7����FA]�P��β���m!!*Q�tdS�ބ[�?���6�l�cH���3�T&;�f�L5�`پE�t��v:O2a��_  �G��vǛ���O�^T��,@ʔã�r=	"���l�k1%��Ĝ��m�ս����̍0_�m��/uu��n��3�������lX'6�(J�۱��ɘر,��C��p�������:�!�Q�����oU_�ggj�^辨��{|�����
k�Ddݔ� ��FU�&��m�]ʹw�P�Eޗtp�����Us�Tig�k�\6ޕ����� �%��#�W�[j@�==����f�q����C�si|�ÿu]��T�H��N�R!9�M�;\�T�@^
�M^_���Xxs�V&��Nj�',�%�g��k.rĎ<��-�����6�9idL�;v�|�]V�y��E^��v�*��M�}ѧ�Grj��)�p���**\՗��7��%O1��ѱ�l{-�w����8������Qs���֝i��)+ڙ�@�L1���������v�[e]^^VN��Z�(ŵe��we���]�Y���n�<0Mt�`i�y}�׈7�K�c*�uytm9N��9��2ni�;��`�`ɾ:y���h��Ͷ��xP������d-6F�S�����1�
G��/B& �N��;������z
`ji���E-�B���#��p�`AFW�<�V�݄B[���7RL�-����,i~�J�Ϗ		��Dm�6Z��R�����A�Ga���hS�8�O���@����^��ٟ�ڮ$)T%ڱ�8����_��<�\�4������t��j�����2՜�ǏOI��^�F�m?" �x ��&�W���9�E+ֻ[	�2��ϩ�1��#B�G��?>`�j���U ��m��A��F��ΰ;N�,*�*���yt��N�V�Ij:�ҡ��H������d�D��%�'�3��w���tH���#�� �ϱ'���鄢D�Q���9����������y"��X܇W�δ	�ߩ�b2r�â�=�nE�ݻ8�Ih8[�ps-6����C|�;J�9�ER-�	[�����9�e���0�������Y{¹�I����Ծz��gd������r=��r/%�,4pU�y+:�O�*�:� ��yǞ<R���e΃W�4&��&��fS�Z�Lc���.Z�@A>�y��N�,$�z�#'���~�<�IzAv}pq�)a7]:#k<˚W���h}� �g~��d���zCr�D�Q���;{�]�z��3��[��T���q]�}�m����/z�91+=U'���C�%y�uv�c��s[�����u0���3=g)]��٠��$�0�������Ij���*�H6-®+:6jVq獗�L�DV-�tX�[	Oq�-D TY)�O8+ngÀ��	1W�t�P�8P�5�i���q/�����Qj/�jY~��Ըq�w,2������~��.�W^�;C���g�j.�p� ��bH�V�qk(y�艍k����bN�W���7(�EIO{Z}*�IaC$bH���9k'�զe��kx��+3����z�DtFe�}7�,)*��q����|2�:�X���œ�����]Yg�^{���e�0 �U��a� �i�l����%���W$o*��PEKe���3�h��I��eo"f��m\.��Iڸ�i*�
��D0m�/q�h����&�%�N�O�`����JfJ��Y^w�����Z���@OJ������
��t��{��<�[�����=`ys��:� ��he��d
'�-z�A�/tT��S�D�_�nw��.�X0Ԥ����_^�������\�gbzY�����M�w?	,�@���D��`���e�n���=��;�_zm��\�M����4�/�� ?�'�K�M���y|�<u:̕*Oۯ��	�xB� �\�&e���)a&t�B��E�L��۽V��7$PZ�ױp��$[c�Մ���B ��/(��t��gU�V�~<�� ��I�z�F:.�4'u���?��1p\?���W�����E��D^-ܤ�J=Y>o���wt#%s��HV0%Ϭ�Yz�O��uul�l�u��}K�e#<�������wc}�
�j���kCD�1��A�����#��8x`ĝ�a�j�#�x�v@�
u3���T���\@w��n<��~�S��ou�."S�?Qj�$j��:����8���H㔐�t>�<� �珍��9/vpsq8�6댢6\!$�>����4���4��u�����묀�Ofr9�ˆ���q2.�Ľ8�jl�z�-`G�'�4��v~\Cë.�&�	��}�n�]W��~`k�f�î|��f�d�>4���E1OZ����+Z��H?g0���/5�*#gV�!��⧵����[�E��-�pM�
�	!գE�����WH�������/K�=.|:9�]+�7Ҟ}�#ٝ!H�@3�#5�`�o;�<c�w<��sT0J�dU�H;������&���K��HV�<'`�|q���٥\H�l�_~;�=R�M�\�J�G���s��H��0;���V�L���D����=;��)f�=ߪ���+���ɦk�b���阇Xd�����9��1ۄl&�m-�m ��qF�([�gj[�(XHR�d��x�E�k}�Yٶ\�u�y�y�]U�)ԃ4����?s�Lk!�a�7��:$)I�^3�ܩ�%�2���o�!�3�ΈJ�F�/���k���n�}ߣr*ebՒ�N8�v�i�'ِ��SOe#/X�1�Z�3�	�(�Cs� �������L�/���&�� �0����p�[�_�F��6@*�5%������qdǕ�?'r�T�͔ȁ�����A$��<O����%����8��R�JL&Q8q�3�+/�2�\P�
����v�gݖ��0�j��61�d}Y���o�� ~�x׮�"�*x?�m�k�B�(h��?�)�UI�	O���B�q됍p�]%��8*s�M�y譙*�|T5��͠d3��Q'��'֑��m�����~�si_�N��IV�T ����)�	(�Œ��&�%^~�����JSA0\$��Q�E���`��"��\8@�����3%NW�-}����"99Cf祧��aTn�\A~��\�m��	W-��|�,��S�T�7H3����)�MG,����'�*�n�{n^�ueɌ�s�H&r���w��NV�v��!W�٤����*��x��������s���Ц�ҫ��CK���rFh����n��W�WF���0DI���d%+4�[a�˘(���K��eE��.� i�r��a����L@���~tl��MK/p����	�8���Y���AC��g}p"�䶜i���mnr� �|����T2�9��2��	����WZ����ª6��Q���e]��0*���Ր�$��N`+���`��s򰾺ú��T8�6��ިg�I���*�j�YjĹp{S���5���L�{�* �?G�ج�Uo���J�U
|s����L�_t��qNKʉ^�`߃�h�^2�>�����%=����	���sD�o]X�7�r�{ d�uV�C�7��)���^��d0�����7W6��jT*��2F]b��7� �Iށa�^eL����2z�� oٶ1sr�s<@bK�6����_����o���Db����C�i���z��&*۝�������7����^]a�w��[?������R_h�{Q~�l�m�ǝ�7�gx�4/�65B���h�bE��N�^g�Nx'�h�bءu������F�J��z�~O�}��TD���Sپ��%��F�w��Z��֕���Y`�4��7�<�A�5Oqu2,ȩh��3I��8g�5Qr�nF����1a��=ø�E�t4�z�B��}s��V��`|j'W[� \*�	�yZ�i�nᾲUY,�r2�N'"����D�b�+�6�.�b?ϲ�q���.\ƀ�Im�/��@�(L��q�d��iւ�?�P�Q��r�� n{S9�� �B2�N�'a*!��~�[��i��tl��FRL7	G3x%�{d��d� )~�˞�*�̺ᾄ��Ƿt��v�G.+%�ܒ�_���'�	ĳ=N۵ծl�/F�G�wV�V���(Q�(�Y�\���CJf�k)�7_<��#��;�8���+8�%,�F�k�T�9�7�$�g 蔉�^�B{��Gt�C\���������X���\��7U�5�/��`�hݫ��̪4�� ����x����t�.Юb3���1(E�5�$U�J���yR|�ά��1_:q�Nw�>]��P*�Vן:����D#܏��摿_w��6�Nqg�sm"�N�.^$+��M(9Q��_>x�p��p��'5t���WK\�ŔP����}�)yM���Nu���k�u��$�d���&�$�2PL�>o_�f�7���1�ň�?@x�RH�	OWh߼h���Z����:��U|&K(R���c���˪�����/��A��w�ǤbW�m���)�EU4f�6�&�����o3����q<�" &"���
@+9[Č��]ų�Wٗ�:־75s=�o��\��%\����W&�>4O{���v~M{���֥%䫓e�ҕֿ ��hE�חt;J4_��2)��\��ߕ�l�#�vd�l�z��KN���-�| ^
��`b��P��3A�T��@34�-Sdu$�����Fr�#��~A�`���qB@�)�u7�x���"�����w�8)ƵŲ�ˍ�D��8���AɄ)�Y<�>��X��,ݻ)�mwt��=�d�l�P�h_�U��� �Z�-R~�*�P{Fm�1�9fx�Ȥ�׺�����k��pt�L��tx���b���#���º	�9� 2�d���h�#����V\6$y4 X_��l���g.H������u���y.N��vw�Hԅ���R¸`��*��}����������MQ	�I��Hi�;C9:V��������WX͵�V`˺���@�7I��3�ڍ+�#�,1�;�$]�a��w��O������|T�lE�噲�4������g�Nhs+�B`����.l�`"�Ph��V�|DBk��V�^+�[&�U�����>���(�t�P��gn�ɛ�^cd1UF�u�yoU�b����w�Էl�-��q7>
-��������kWv��4��ܷ�;�h�#�C-�8Žo�:�e�lt*���Ԁ8�ˮ��옮"ړ�ԅN^E�_��տk?��J�S,4�oah���F�*�(�[��<��	�֋��ĝ�����. Ģ���<˗mjo��b����.�a�Qw��X�6UlC���}BwuqC�Y�����}2�By\q�������B/�>aϝ����b'I?[�p�M��S�:ن#��8�F�=������^�����޹K�{�d܄ǐ�n��oDZ�{<�UE��J��p��O��ӛN�=�~�A��}�U]�V(���vS�>&A>Ieč����:̒�ĩ}p��������C.'�����-�Q�)Lw7�t�A}"H�AB"W�"l��R�^�9���B�n�����F�jv-c 	�.@7�*�H�g�E�*�5:�����]_�H���4Ԓ��H����).z�)|c=������F�&�x�S������R�.sa��̆�$�^��=O#�@�h��o��9+_5�ӡ�:7��RG����:R����yJb��#ݢnSa��xc��	2�U}�$,b9ҽФ��s��.'���^H�1����̭oU$����]���7�|�_���e ;��4�U��H6<Ȣ}����s)�h�)��dh����!�$%�|�A�[��uu�M����'�8%D��(ȸ>I^CvކO����c<Q�`���a�ķ��\�3s����dP�0��د�ˁ�0R�ln4�p[C��.5��ߣ�ϙ��,�w��𘫁�$�u/��by�(����,�RZ�i"4���	�:�v�.om�V��@�¢����.|h�Y���J��<���y+���c�++��%iV_�3�=��M����,�Z�0(|P�gu�h�/�&	��������_��h�r.��`Pr"�y*l�7�7��sͬȁ|�Z�$�JB��5cG�}T|ФqCh��J2��z�;V�Pۦ���%�����{��PԄ[�B5߀��D�����Ք]���
��?Z�\��K��v�̃���wi�|O[K�D�J^�Y��
�%�Ɠ�6��_ U�"��v
T��FM_��p�u����3�_Ј�.|Dʱn�:̌����T���y�E����m�0ĺFy�]�r&_60�*��d����״Q)�+�x��c ��(�b�N=�F,��
�~��GlINʄ��ӈ.�7�O1���J���q$�Ee�g�<�J��׀D:`�VPH�֓�2,�3���~tعT�Պ���t��'�*����j�N��ӻ����>��0�7�h������,o��_�!�,r>R�|#R߷=d��(�Nu�5P$,���l�R�W~��x��|���ߗ˸@�����-��">\���m�Mih���.�̻�Z�5~�ÙEm{)��2����xwU#j�v��T�_�����qB�R!����S_����6"�A�,j��Y�>���Ӣ��*���_!��k+w����x�c:�a�F�|�RK�p_F�^���,��"��زG[	��Gu��'A�+!�Œ%�=V�B��9s�Z���˫�>T��X׿LY�G-��~I_aCM"2=&6��'�Y��̳�Y�9K['g�)�����!:)�_��w2�v�rwn���
uN��)�6
H�]b��N/۸Sw͎`]|ض,@�OhD��9��NPSi編�SI���kϥ���Ʒ�j�ć[�[h����e&�u�e���*�n�b�s��Z�j_ej�}n����D�~��a'�<b�'u�˸��\�ߓ�ꓬ9])nL�0X�B�E�LC$���x.�Rooѿ� ?�$m}�VN1w�X�W}�g�7R�iVA=Y�2?k����\�&h�����SA�U~�|-���$EN�p�qTi�z���0e��e�K:8���a�X��,�2�gu_?��aSO�<���gwK���n��R8T~l��Q�QSh����-�6��Nk�T'P��^�uq�W2�/����\52K��� w��|���s)����jy'��Ev]oAT���^OP�7���!&�c�g�|��PxLF��O����ବ�٣-[`�r�N�\f��t L�~R���w�$����9Q��h��[�~B�Wg�D��G����t)B��w��d��_��1�и	M��pf91�B��'D�I��T�3���z�r�$P���:[�V�D��Pmz3�<�4C8���=��ٗ�EW����(�l{�6χ��a1̙�M�.�<�W�����G/�P��-[f�J��_�ͼ��yZ�����}I�L�S�2;K+�����8S�p%�S8�g��ͦ��M���H�֒aYJ�fW���Z��ysR�J�a`O0�Y2@���z��`�������s��V)�Q�_��E�&�J6V�m�����-5��I�?���D�Kx���瘮�03�?��m(��q�HN��?�X����z/�혙;�jq"*^�|VL���]J���N:4��**4_����F`<�>�ːF2�}YVg��9,(��Tbf���T�R��ݲM����5s7�stL^�(GW	)��E>r�C�Q�1�ȝ��D7BB:=��Q���S�.mT=Z���O��_�;�j�묂��ftY���&�_g~�vA�M�pD����M5}�M���>X�$ݿ��w,���%��)�ˎt� q��d{qi;������$,ݍ�H�+��Fj�VCr^ ��Fd�#�y��{��c���l�T0M8w��MY������c�Ȉ?��{ї�~��T��rZW�?������*���j ����*~x	��c�r��;�� +N�&.|V�r�A�4'�V��ʲ�J��{���0���^L{ۭ�5�.�k�'+yu�ᝬF���+���Z�U�G�W���o��6!�y�ÄT'���ٝ����uAgZ�Qm����/�<��yL��I�|�V�Ch�b\̊�ےK��	� %�#���[��W��h���9܁Nm
b/	�<'�����xP��Ϭ�}��]�ø%���w�|��ͳ�*S�b�6ߝ_��+��C�9��J���ܒ�g�<	��91W�}�_{R�|�����O�t�����5��Iח��jH^Q��<��
S۶�g���m�wx���~���t���c�b�|�vJ��vH���!��Ǝ�������c��/��t ���مw��j���cu��N�����ٟ��s��g��j��������-�]�a��~Bd�a���&���\�AR{���hٌ�v��Ҫ�c�r���e).������@���������i#'E@Y��z[C+��0+�H�o�I����7���Rd멃|��@1G�/$>=A��Sx��5(^Q���
5�A����Z��:i�EZ�]��<UD��_o�X�������ڠ Mx�s9n}L�no.�2�!<�RF�4�5,��h���7x�dU�>�O�(��
��>D���r��=1W �S⁌�������/����Y��A����,���m�*�)��H�2HP�b�j�5}�t�x��#�7>���i?��4Xmw�j�=K.L����X������0܎������y��A���l|Ν�_�n��l���w*��֛K<�5��@U|6�%�sFGy`(��/^Ճ���mYA��������I��T�T���E5����A��������I0�ug�[�ѕ"�	M�M���R���BH��r������>�3{��r9��r~T/��`?�;�^б��M]��:
��n�`7*+�D�Y���W�̇-g>~f��.�[V��|���؝@�O�2�8?'����d*pK�/��Mݭ�7+6|������JR�88�ӗ߃��!�����K*+��H��&Ytݴ}�72�RO:k�D���+Rе0Ţ,.�8��c.o��b�YC�eqX�`���l	V/��z�d��P3іiQ���tһ������Hjv�S^<� .`�H�[2�����2e�$�sCSL���5����5@��p�X�����u�-�w��dYL�̗���q�_�?I���4�(���[���ތ8�����N�ܫ�iGbB���W_r�$�\�P��K�������Һ�7� ���/jV�~��������{rgu٬�ǩ�6�V5�Մ��r8+��jRA-��
��ϑ��K�	!��ZoV��iΛg�(h� 0Kt�^�Ĥ c����M�f����`a,�X��;�L�R�q=y3H|LG���Rs](ZV�2�������߶���$�<UƠƋ��A@���\�i�AE��U���^6��jaz��j/��"໩W���§���R�d=�̯�'K��F�+b��a��U=_b�b[:�L���m����ZLN�3�p���O���-�0������`�� ��9�RQZ�,@@�o�L��֏Z�9nz�t�8lϪ�XSFL�\�\۲�WDK0g��;���6�{$�r]�������M��B�q�Y����t�Bj�mW�x��l�RnS�#rQ4I�'�j������=�֬�����1UEewqC0/_�ƮW�ͳL����]���!W2.��UG���x9Ժ���D5_NeδTɉ?/��vw~]���'�܆����И,��p�-��$(]���?�j����;t���Ʈ��<T�
�9X���)j��.�2?�$ӗ{ �*�c�a�������Re���5�%��jl��D>w�F`=v��#��O�!g�ie�9�0fgtf^��d��<^$è�K��~�wn��}M��ʁ��#�cdJT$�˚ox�}x;���>z�3�z*u\	�ʾ$���'U�ڨEL{F�E�[��`h�mo�ȶ�<�H� �m����^)ز��F!,t�| [Hg/���s=�=�����4Xٙ(�DjL�)� )��� z���w2�p_A��3�A�@��Ň��Q��#o��5��Ϛ毱�˂l
�;D���3�)�Qu����j�������ײ�j�3Q@���D_�y��}��|��K�B��U�w&�6����x�Ũ^����>^t������\B�lV��5SRL(���!C6j�2	��⌸Yr.�9]����iH���7��D������#�E6X1�����EP<@X��I�ɥ��Tc�l2>��{��Ae�}�����M�z���v��:�P�X�G�rL��=�WdG!����0��dD�˩v�A��"0��]*�_�������m��GYG����`;���ߵ{z\'��!<*�	�3V.F�tN�T�������V$vr�!"&5��EH��~CE���
r��&BC"[تEM����3�֧|$M1�R�Bh��\��� N�ʹqM�-{��`�q��}��$������=S��������� ���L �vWB�hYk��R��K���2������iG]�4�������<�iL���������E�?
��Z��W�/�>�T�Y��W�B��_¦���N
���B-��U�ށ��򆃺�+�<�~h�Rc.-*�>�y��Ͽ��Zb������V{�t>A�
�+·��OǤBil����k��� �tk�W�ͦv�1dҡ=Tf��Z�G���a�p���Ie!���U�H�� #$�:�rs	k�����z��R�6�� ��]]!G{ev���z���uuB�.��!"��=;�ѿP���� p��&�K���|�ݣ�
1��ʸ�  ���cb@SE=C�ݫ�F{����i$�G��c{�oZ�'&��}�i�
�U�t��yy��V��2-m����7RJCT��x����)G�tsg���c]�­O��Kh�G�b"�Gz�g�+J�at��e�����eȻ�vn��5G��B,�6�v���<�DMeX�Ym()a����Nf)GL�H8"x߶�>���XmI���W8�2���s����]_%�3o+��"Ow�#�y�
�*yˊ@(�d�NOߍ��wcO���fc��l$��2j���������:Vv���W�k*Qju�������uF�QuآTci��R��1���Y�9�3F[�����PF���N�� �O�V�z����g��`9i�&����2)���V��� �7��89�b���|��d�㏠Y��s�W�HG�D��A�d���X�N&4�Eg�9�a�_{���C���5H"9��@���(U_inZ��3���1�'��{�Q&9THs���a-��Ag��&WaT���z��m�ߟdL�`��%V�d-7�1��V���~��p������l�N!��l��e�p�n����J�Ω?3���D�uqQ�a��٪�hǇV ��.��;eɑJ���j����t��E2���Z�IY���33����g�����4-5\�z�6���<���Q�H$��0V�`/a����b2��n��k���I��qG��U�g�/p�|Ө�PV�4�L纘���/���ixZ=ra:�\-��%�ݸ��W��g/	;��D�]
D+&6��{�G.�nE�z%jmu�f��$仴������0�D�Aa�"�o
��������9]��P���ǩH�(�ĳ~\��2�b���<8/}i���* ��A�X�j.���U����*+f��gw�$vc�x��̙�2���Ѻ���ke�u��1S�7����l��^�+��}��h���1�_�+|�ǫvcq��[�oXw]��N����M��z���4e��`�,]�����Bz�E��������}�<�O�i5s�Q5�gC�_2H��B�o&Ĝ�m��<}�����GJ�γ'�����o'��T�e���*f*$
j��qhD5����~T����������pھ�7�����.��_.�j�=�)d�(w��d@٩��5|�A�\�N=�Ѯ1�/��GHEn���21� m~i~s4z��"?fRO�Rc���U�,=3��fӸ{X	(6h�9�qL=yȳ���Og��9���гN4�QK�D��U� �;�UV�|�|@!��,�Ӿ+�Gqw�<SW.^U���Ⱥ��j�d���d�x�	{������G����3�f:.�8<��s�JQEg�	��w�[�S�l�eh��ͥ�55�nm��E�M�l��O��8}�)�px��@��au���G��4x���]������ǫf�O|:%��p9��swPE濸�,B"m�˩8���5�W���<#^��^�	��Q*Bܶ��lu�J�A/t�s�����m���;�������T�FD��M����֜	:;���k�e�I�#զe͚��2S2��3%�K����=:�n������h�vb�)s���ԕN7��dU�i�)n���D^6i�a��e��X���t�u������#����Q�hL<�+|��ɝt��P�^���_e�Y��w�v��T2��e��虫���eF�>�PX*:a���EE�D����o�+��rh�U��Ģ��1�z�wlO����mH�U�
2R��}<V�yc/���:�N�':�n����
��	�@X�6��>>Mމ�Y�_r���F*�-��8��\c�G��I
�%D�}�RdnV]Wίkc�N~�y%�d/��j=Y'X�)�t'�|�!v���y��A�%��� ���Du%)�^#*zX�rI�p\��zL�MwnC�wZ�E�K�>����P����D�h2��m$K��j^Ds��B9$�X@t���HN �6#��Y���O.�t�gH2�D�%;�U4A~*s�)����
�m+ ִ<�A��%q��2E�y\IU�[�Ȏ�%v\q)9?<6Ιo~���(��4�t�����:g��;"<���u�}P[h5������ژ?x�_�RE���S?��3�se��u�oD�F����+�=�oq����"YJ������DP��D�-�Vm��Gښ�h��s�}��w�~#�P�u�l��2H���!#���j#���QM�*�;�evɣ��b�E7�%�S#��[��T��t�;���&��gZ>�#�9�|n�����R��\�>$�Ʈ�'H|��4c_��E�M��b��J�H��~s��8+��M���m��	z�3�>t����1a���/c���2B�I{+; ����!y�L�D��l������r@����?��Bl	�k���^��0�._�����[Q��m:#�8�g���m�>��l�$��O�Z��.r���+Rx��+wC����M�R@D�O�yQ����i�f�&|;�SzW�N�"��+Voy��-�Bz��Z���X�Aa�����ݸ��D��el4��)�tX,QI���V�T�/^7��M��	=����S?�h�r����2���|��M��1�K��/Mn�r���ྌk���_��pCx���5���yNgÔ}�����fqLGa6&�5���s��|�K#>�MA�-
�7J����RXYi	�@Z(~&L4�j#�n�+�T\��<�/����G3��z��%S��U�87�w�M�ܑ���z�l];�I��K
���fMeVHKFp9�qD�Nbȳ=&���[�h�����mh��$�k�ݖ��ߨV �$�<��Ќ+�m� m�n��[���3zG>�H��Ʊ���D�10�V���a*�LDO�baq�S �D����^���Xd�5 �\#�O�\ʠ��.CWr��R
�VvG��B��!|���8}��K�]����i�3Z�5=���⭩�񈿃�4G��H�������D��pz#\4�[3�'5�X!嵚�N/֔_\�_9�"չQq���~�W��	�ʬ��Lܯ|�upԇ�6�kJ�l?{��Zv�������ϥ1�)�%�Ŧ���)պ53�7�ʞ��l��mV��I����J��6_�VJr�U]�O6!���,������D8�WR�E�پ��8��F]�����Z!�1�s�[�|�ā�&� ���疁�CK<��GA	lO!�l������]T���af�W�:��26��I���\��8� �fL��/�Y1��Ğ����{�ܫ�A��æ)^�	6�E��/�I��L� �1NBq�nxo���p
�Zt�'>�d�|Z�i���l�˵�o~8z���jo�Ux�����(;ӊ�[b\,J�'�����㌷�^�'��f+*s���^�"��6+���i�}߱�����[ɡO`��J �`���p``�j���I���l����Z�^�H�1¿�μ���R0O���2��q6������tM߫/�D��y�0C"K�$�&l��L�����������屮1��h_��ZU=���&B����UӏYI��σR�1�?u���PA��gf�	�������`9��H��DT���a��[�T�f���&�W�ĺr��YG�m�2��B��x�uc��
��-C�7�Nבɼ���gm�暟7U�%ݺ�y3r��nu-G9��%XJ���zg�m����~6ٲ}"�\���w��H���B ���6�mk5{�M&u���K1n�6�+`�q]kF谐 S H�B��HLa�
8<�����׌�$Dc�����g<l�b���麪E;��W�w����P��>��-��"���\4z˒���T��ϟ���̷cnu��@�6_��ҷ�}�b#s*n��yY~����3g:t3�G,�hm����t�F�r@j�-�
wu�"�0�t����pl�.��mu���a�J!����g����)0Ȝ~[^�O=P�4��u��#-�����k�q6DW��4�����<���m����C�Ek�E���9�t���j�]�Q�gU�c���9]n�f]#;��8����?�V�2���Ҿ=�v�t[�w k�d>���O��+Q��*W�&�1�>��;����DiSʸ�#%􉖛�K@��'���=�ݒ��W���
�}�QO���fLmڧ��s+B�U�AQí�q�p��:��}���G��+���"w�ߣ���JF:��MVc۾ӃU���>P�hй1+�Z����
vy�����k�z�qз�WC�F�z�G��aÊ�!�x�hZ���y\�g*����9�o��0���[�&�dy�����8O,�Y�c[�vR8b�+)�S�B0{��Qx��qJm��!�F� �|W`>~h����AN�q\Z�%c����F���㏜���6SaϐQ�#;�Y��Wlq�V�����2^��=��#;��?\�sf�����q.��;��Yd��b�����|���L�c͢�����c9P$��Jg���,\�����4FVv�cx�&���d�߶)k����?�66뚝��Ɍ(r��o��b��wɐ9v)�(��拂����\'�p�$���#�R�B��W��o̫f��_��Șd�
Z�P�w���@��;���$c.?rB?[�-`��7����}���g�:'?��h�
��<���h�B~�ec_t���Ē�8�s�Y0�@ҋ���Ŕ�Bv��XX��,%��U@�����W�NMۙ���a�<sŴ������-4L0��+�Ԣh[�[^x ��x�ïo�}���������|����~j�/DY�;�����h|��[�XY��5Χcc��}�e9�#�~�)����b���v�.����D��*t�=��a:��T�ZGq�w�pÄ�^w�ND8l�d��:�]*}��"6Q�iQ�v��v�$Fg�hR�j��lSZD�Fќ����>�:�!��+j$܃�~��WO��R�3�O��_C�E�?���.����9��&ٶ�o[i�p;��%�hΚKp�Z��x£� C����%�-ی׫��uϭ�^����^�3@��������ߺv�
XN����ޯ	��'6�[�0Ĉ�����,=�t����4�Glw�ڱP�q~	��ػD��q�$k�'h4�''X�a {Fn��	�e���栂���,��FX9;�[E���`��j�ѨH=�.��ɉ�[Vd���)�{	�j�G��q�'����)n%��ʺ����/�3H)��j=���ִ;��99$_ܤL�ks5�&��X��o���hۤ!mTgܱ�ys��6
n��6Ӫ��ajƵ]�v��P��"E���m�X��"A�B\�M��=ѯJ�����#��N%c �Fh������2Ϧg���E�w�x9x?cƱ��z"�������ʟ�zË�B1k2s�db��9c�����d���r�8�4%C\^�_.�5��]a"��� <��)�<���<�N���[�va7���k�{$#�X�펹H��2�1�{�xl��}R[�m�u�������\�MH�6�l�'a��1mju��M�<�Ms.��w�B2*MV��3�y6K3 G7�`3
��*|.xt��*���Э�5�U��VXf�(����"��:��xd%d��T6��GM�Q�q�����j�줔c��|Ӄ��ā�ܼ�ya�yo�����Q�O�J		��)��/v�С'Odkߕ���˜��@�mN���Aʬ��dr��D?��0��+;�v�$4:��� �O�d�OЪ?�q#�u���K�D&�T��)�I<��ēSH�{'�� -#�:E�4��#�я�[)���%���${+���I��b��Ҏ;����J�P�7A�&�}��K�"�Rdr��x[]O�W�d̛���j���K� �S��8ʼ�����o�
��olŉ<�Ah���.gΞ�?u%Ӑ��r��R-!�]�]Ӫ�j��N��LP��p��=w1�u�~t�]'Wv��,�:��Q?j���@ݝ�ӿ�Ec�\�P]m��&ڄ:Ϣ�8��u0*�i'��:�M��/��x�XJ�	VS����Q4�q3dٮ����]��� )��ʤ�iL��T�C�]-��~�0�	�
�{ų�~u�5���C#���C��$���;s�!��:��ej"�@��@�/��R�'(�Ǽ,gU0^<D~��j��k����FJ�n� K�g��G��Q_����'��^��M���QQ� ��^)��5C�;t)��G�T4zn:R��zIn��J���,!3��H���5x෱@n6'��谇u�>)��5S"������ �`��, ����S��=I�\�KG�Nv��/�9ո�2١23o����0S���o����`�D�;�H���N;�z��n4Fc��鹷{k=׼q+�c�`��7��'*�Mߩ&�h��֭�\�����R�pj�b./M�yȚR�!)��w���|f|�a�8n�I~܏rWh�W:8�L�{��]��W� ��*��X_*Ѩ�a������{@�%�{M�LBt+`��~��Jɕ��%%��|>0��m��wi��de˯����Sޑ��7�k�����B�)�mjU6�_ǖ�1�)�"�Eɇ�&/[hL�@�������suo}Sz��=��i*�Eo�@��T|���x��k
��w�j���X׷�n.ui������:a��ܙ�Ob�$��9�&��"�d�5����D;zC]%:���m��xF��\�����}����nA9�鎵|	F瘯O��zZ|��c>$�n�UN�����==����g��P���oQF�����o3$�jzQ}�5����0d5>i�{���Ut?��nw0�Q�X&�L׽&�d�R���.�6`�Ɇy��箳����Л����d]���e�.Z����(�XR��/V�4�8lR�A�b(��4�#���v'�Huɤ�m�r(��p��������Rg�˲o�����3����A���O#��� 7���b��pWTt⠺�@�z��@�u�9���3�*��!�oek�=3�{�b!������Uӯ^���|c��,t����P`�c_rI�1�r���"ݤ�$�}˰Р[+��>��Auj���{3�P��[1:�$8�c_Q��[溢�ʖ�IvQ3d7j�W@�Hp~��}$�}�l�]�f�m��~�n[��! А������B����4Wy���^$�y���J�ru0��Pv���U�����]�1TC;�`G/�RLL,��a$�C\mI��O[�抆�K�S��&��}+��Љ��OY�T� �XC���Fe�I�n>H4�i�x�dЈ����c|�7���O��B�%H(��&���#iKM}-��/ ��i�ˈ�6D�?�uw��#��L1�5��ߛAڹ�tZ�:�C?��:>p��̀{��8��U%�����4�\�u~2��
�fV�����7��n��@F*A?�s�z[�7:ɽ:?�8���U�l\V~��Ȍ���l@��4�㖖,:=�?�!���������=-��&v7]_���L�̯�� W���`�)���!E<p�;ݪ5G8�d��yuK�1 ��g<B����S7�$��[�=� ��R��{K@mʃwl�V}���~:r39��oܡL��=:?�1,�p��ѕ���x~��8�"@�2�6SO}+�}����r�;�D�B�v6=�O9�	��	���Z��A�߯e���I��;�s5�,�t��u�y3��B���cp���(|��*k��%K���t��}�y�y/��Em�����j�F-�]�O�����C%z	�Ƶ���v���!�J���C��H<�X�k��]�q�:e��0Ԟ?t	F[~#�����d����Ӄm;7��v;�	Z_)e0vI�ˀN��2'5e-m�Aϒ}��A��q*س �H�������EF�X�|�	�Y�*CJ���7�**�<Qav���zCo��[�o��id����:�F�ϵh��˟UY�����Z�D��� �!B�s��6"����/+��F�s����zI�V���.���n��W!dYN���K����L���iͮ�
(u*`)����d�֐�*zX��X�+x$2�J )�j�\']�^������8���u)���l������ ����w�F��7��d�qY��
���j|8O`~��6@��	�k[��a��F 	�uY�ҡ{0�[�N�:�������t��CY�6�	͜[^lz&`���e��x���6Z=�d�ݍ�{��գ�o6��`pn��^�w����F, ��V����e,���~�o�R�d0��l}�a�
�%�����]\*ۅ���}YD��GF=��;b���O�jb�8ܜ��
G]]l�r�o�͹���ܬ��Vj�qZA���ɵ� ����u��8��oᷦ��S�&�%�'iBHX7M���w2��4��@r'���]�W��j���qA����z@�1��+��!�����F��x���7�Ӏ!Qe��y'�r������.�S�>���e�Դ}{
D��IP�͈�#��D���L�LlrX����Yʔ��:r����X�*�7�i�EП�p.�T�H���	Wa�u�/ߢ���_�G�p���}Lj�p���~�>	^����z\~,��M���/S���߼g^Da�,�zh�#̒4�P�N�6���nG-Y}����- XI�hFΆW>�)�s~5E�{�N������Nv��W�*����M1wP�Q�dͅ�����E>��y�
�,��y���z0�M�E+�QY�F��(z��U,� 8���a��?��v�gi~p]�ѽB��I]8'-T�F��Mb5�<��n��G~�"b�4����׼څs���s�TE]^�dG���Tt\^~{�jb��>������b�d4��DS�xTS�q���P��%#������Cb7����d�J}7m*��A�:5d۬�D�=y���4�b�@� / ]�H���Y�M{v�*��o�]�\K��[�dV�k�_I������<�����h�c��G��|a��_��t���q�nO��9�4��s���(P��
�N��]DJ�+��avq*X��a:��6��۹x�Rw7(�aE�3�~@?�*���O��˅'�T����]rLf�	���Z������Kd8����k֢�ʎϜ���w#�Zo/s(�oW�_�7�u��s�j� �����O`�t��<-�B�N��$P����d	��$y��l]*e����8�c�����@�����)���x;�C�eAٱk�^22�@e�Li��3�o�V)�z6��>[���8���<�k/~նӿR؂|��:�D��]����7�/
��ﺜ0͢�x$Sc�|&�u&R��Tm��������X�����Q3�4'�}I�q����2 �$�M�Bpޝ������4nL^#�\8���7�3�Uښ�K�K��ր-��ͮS��!Re'�ʬ&��7:[�Ggҋ'3��X���C0��ߴ���֫ƛ�h붊�aw�'B��.l�]lYw�3�#���9Ay��%���Z*2���"'M����E�'F���3��Ä�.R�.�ʪ���eMHz�����'_cd���ڻ�;�Zq~cR�u��U�5�Bz�V^�/X`\�̡����XN����*�H�s�Ce3�+�X.2z����:�3Q	ߌй _A��L���ʚ���c] �Zr� �� #�YÂ�Z����s���!U�; ���Ys?sW	�壤(zt�-m�:t�ۅɍ�ꃍ����5A-S��
z����C~�o����]���J�"fb6�if�{>Rb}'��C|dJE;Q2n��n�'���t��2C���{�:ׄ}ރ�Y����L�;.�ID9���k�V�a�GzLp��E0��j�B�vN[c���x�LL9�`�\�R�w�ێj��߱�}]�˜������1U�}�x��k��hg�,�C����p�?c[s�}vc��0�����t�����{�oQ���0��e�c9�|jк��
��B�Ž�u�l��5'�-p�Yᣈw��82c o�eK�J��@yn�:��n�5��{c�O���'_��f`M2��}��&N�YZ�0������S�B�O0}��61��7�� ����!����B,{yI�#��d�v�V�w�N�%�r�s���0}�,xH}r���V/4)|U�#�b})��釔�e��z7,	�_O���-��1Ձ�X��=ׁ!F�mƛ�Mp�[)[K?64N�~|q��
ֹ��A�ͱ	�ҡLY���o|o���̆�6}�Z
Q#���鿲��H��	��4
��� �vr��|�F϶��0!��7f&�e�uͨ,�VtM���r�
�c��]���;jG�Q�AMH��k&�F��o+��(^��@�P���c ��8**`�JV2���tW����f��aa���!F��h'�6GCFoxq[/T�I�$o׺|P��9q�_	�ܷ���LWgPdK<2(��J�)+��/������[��~z�\F��x
�Ũ*��P<��O���A8�œ���|_�ш�e���:��{>��y�{@4B����`��տ��^eĒ�[+��9ph���_}�?3Y?�0��tiި�� y_���2u���/�W&�u:ee"鹜r����E���:妜3��xlT��*Ƽko����r9��+����-�n�WXy"�z�q���e��_D��B��iu��:L�z[i��-��[Cg@#V�>���d���6I��Z)�]^��_������� �Mm�����l�ɋ��� z�V��P`���ڏ�c4��i/#��vZ�нf�n=��B��<��3���}`#����I�=OB\|��*��'������E�*x-��I���J[��cU[��,�U��'�nL |�#Dx"��N�.x �{0g1�{����Oş�@p�6��\m?�mU��N�ز'�F+�C^7��'������f?��YV����M�	i�{l�[���t�����B���!RWf����J�������˼��k����Ѝ@�s�a���;�ex	>���1��n�	�8�)q�'����.@��v	���p<h'N�`��F����A��N�Y��#p�O0�Sr���^�3�+|�d]���eT�>Vj��q�v('~ɜ�U� �dj|{���O�z��K>��M?D���z�GZ�a;��0���0{F88�W � ~�W/󩓡��� �$�j��K"4�fQ״3P�pFp:t�,��"V��a1j��Ej/�Ώ�&�i�֚���ܝ�����E؍��Vq��C4�9��ֹ�w���w�2 ;k?��Y�'M��ߢ`�u�����s�r����*
`��]*��ia��[y�lx�߻l���9i���qFݎ�2��GT����}�j��	��7�Un�'k�/��/>:��,Nr�On_���6�~��@�	Z\ۉYp$���jw���q���su�<�%������Ҩ� �:��$�=Uz?�b5��d!���9��MԆE��cmaз���p�F��-�[�������$�ܨ3ȭ*�[=6:EmT�pu��QZ}�Ki�y4���ͅ
�c�L��<�\3�!}�_{8�U�|N�B�[o��<X&4�0"<������������Y����0�m��!(lr 	�i�ڻ�r�	Mс��b�}lg{��) �ε��λGV][b%	��Z�ղ��.�a՟�S"�M�VY�����*J�X�k�ЃeU��{o�O��TZ�^���bn���$��%i�:hl<�zDz��Ť�u��lf���=�cŲ ��/���#</��T�G�M��H��ORPI�.��S��-(�a��d��չ�܌�NL��<���K��^�OI�i���a�j��SڨLYV%���dq$x�}~q�g�^8�Q��d��:��r�  ^Y��W\�$0�B�cc��W�qCy�zh��u�檚o[K����#X7_�KHu)!��3��D��ǌI���_���֘����Y	�nm��7�v�Ԩ⥇yac�N;Ex�T��l�K�tC�Y`o�}:դޚ�Ft�ބ�%�n��	+\��tzC��>��/���u���H@�Ŧ��2 �����j
����E��wH�CK[=��F�l��T���Ο����kg��F���������2�y�����:������h���Ǫ2��d+�|���A��>X�F�%cX�M����3���t%���c.���o�^X�H6�D�OUB�1X����%�eu>�}ro�x�N
O�睨-���V+�R
p����ϗ{#>Uk�uxE!�HG�g����Zk�E"�1�;q܆��U\	�@�H`)��xv�|A˲7>q ��5Ӌ��	3� zb4��ߩmo퓁0-�|��G{�6l�vaY��n��4��n�s��<oU��,]�
O�����@S��wrh�W;'�H��K��n=ú齲�F8!�#o�$���H�(w��N%y�>�HO�S��o����O����n�T���I�RUX0�ֽLs�:��q�G��Q̾wh��!xj'�l�|�ƥlpp-P�>+�f3��/��|��]�5�F ��^vS�W�ԋ�7L�_��(���Ʀy���4YO�4t� a���ޱCS��^��Ȁi��>��8�����џ�������5
:>���vW��A���TEx�^���`V�n� ���x��8l��G���Q6N�m_��As�i�[1��ph�-c6����|&׭�!��>؁Tf�I}��uF�
tҬz����4�����T^�Y@QN֧+�0�~�F�M��|��q����1Զ�H�ծ�}؞U�S�p�w����'O:=��m�)��Px �L�k&tɁL���Q�D�V Zr��������T�\����0]U�Y�C}�QL՚�Ե����{��J�I�w�zN4�]�� �^��ű����tE9>�ڑ~����!�z���~�U�,.����~��c�m�-jv����#`w<��b~7(����X�nnb���̒�nq.����WX�K�fn6_co����QQ��g���_h�5���!)��}"ţ�̾R[�+�q�Wg��,	���@C&�O�uJ�^vK��"�a�{���Y9/�422�	���Ս�������K��D�0h���YsQ�t��E7ʀI<��kH�lj@�" ^�.GmB"3=�p㖗 ���y�Ԩ��"��O���Dq�����Jo��7�3���Kq7�g�!z[��pսr2�C�%����EQ�xY�E���'0�i~�	ěn]���?��m�s䂢ȡc9﵈��c��C6h�n��q`ɚE�Q���;�*3$֚k
8P�DRAaNC��Dw�=3Hd ��Tv�ze���Z~$Ux��J���/�bb�m��O���w-ړu7�6m�$���� S��W_'��Q�`0�qс���@剥F�M`�^[��+z}U����w��t��Փ� ��8��K�֑v)֢� 
�z�^��7������ ��K�!9%�1�S��_x� �x&����U0U!�?M���~�?v
�K�z1�Am���$P�M�luK5E����+|�����e:��|#�+:i��atE��e�u?0Q�0�a^�K��H��4|��3�]�FڦA�:�������YQwy�f�f4#����x�kN	e�w����s���4cel�)�v��+mT��$���qa/5�9e_�Ju���%L�@5~��{E��S<�y��,��f��r�!8���S�]"�\t���i���ʔ[���o����M���B����=�q�"0�_���+��mk���k8Y�bLGO3α��Κ4�|�г@�僧���(Mg]��IR�V�;���sw�_�WOu�ے�ZW�!�`B���Nw3	MŇ�[ʓ|�o1�c廠dO�*��$@r��M�/<4j��0������E�U��˭�'�礔�ߤHҼ���!A)T�hU<�o�cߧ�EP:���zw��fP=5`��:�/�j=��!�?���P�߹����0xS�_�x�:�ͼ`|����� �ᅱ%�ɍ�2,�Ӹ�p��.ў͎N�|���:w�;����JW������ǰ��|Wl9��P�z+��V�`C��!�V�t�ˆ,�~�f5T��RfT��=��7u�k�(���K�_��/��(�����������r?j�\'E��5���������@	}jV_G�l�X��'�QwǊ�g~ȃlA�Is���/�$�;£�=\;QYf����|7BT˧/���'�-�GU$���R6���mB������h�����p��%�u֞�@~'6Hd�C�s�"�4ni���*#FP�)Wt�B�Q��,��1�Y�#��&Tgdr\�Ҷ"�/��y��n5��F,o�$� ��������OU�0.�
����;�{��|(dn� �!�-�W����¿���W ��%�:]փ�s�ۥ�,J���
�%%�h��˞n�#_{=<xPf�p07�׷�g�x%��u�@�s���n[���/!e!�hI��7ŘW�LNa��J�ܱ��r��o�"8�� ��IX�&v�z��;yQE4#]嬨�P_�{��?1Y��7�S%����kPC����}��O
�2��> \�����}�D�hm8�O�?����/�ŶM�~0�SI:^���W[��&�Vs�f�4YO��ȹYֆ ��,�^��m#�[�����ߠYPI�ӯ��Z���IN]c5�_^EйP�m��-g����;�L��O��P̪���%U����?H�3�h����a'[��|�;L~�����(e[;B�'���d
2���,�%��U���{��-ja~Ӓ���a�E�[���}2�����"���-����>�Hg$2A_��W��8��p��{���P+����LVzD�*�����X�*36�rG{{ϓ|>5��N���芚5R�'~Q��d����j�a(�ǯ�����T,��Mrs@Q)��#᣸V)O&�:�%/&��.�ߚ��>�t'���re���->iPf�.M�
$���6D��e�~�*�?�7Y|���R<G�V�Z<�5Td�q	5���k�z*h��$��^T�l&FAO�S®i����_�V�*��y_>D�?��\�SQ�oPBC���C�lP��`�E=�����@���#�	SZ������P�/(��#�඄$�M��g̑�'BE�0?��	$��qj�/\��TDcb"�����F����N��I'�ט�o��?��׆7k\��IYw��W����W%Rx��D��|�@#G�v�Bu�T��tr��p���R�yH�{W@y?3��d^���{�?�B I�p�쫼n$��,�5!�U�G������)�c��D����k@�?�koz��^���7�/xa�zS�������P����u�"
Ƶ�?Is�-�`���hڌ�3�z2�o���Լ����Bg�r_ʰ��jA��;<�ۍJи�+�z��� ���!Vi�w���ۆ
� ���D}���i�l�!e�G�F�(u��C���4�ԍ�[lL�^�c�tUl�Qd�� �+��@�"41��<��#T��E�Ӏ0�\F�;~���ܞ�f��-]r#�w�d8��B��q����/2�1�����*��@�"�8�����d�ݖF��g�����n����,	���]>�fj�F&en%�Q��v޴�p��\r���t���q_+�I�C9�ۑ>����}�B*�����;S�4P��Z�2�F�k�N�M������a��Xێw]�k%a����uu�e)��}����||��w�]�y�\,��%p��,gyHe���%��&�ƭ�=��,��>:�:P`�Cn�S��gBt���0�N�<���JX�"a�+�'�p�$�p��L@I�FGf� �(�M��\J_`��xI�uy$+P^������>$AR?6V��ֺ�)�a<r�I��-0��ջ�0(� �g͕I�?��,��ZW�� ��oy��M*�[<d���ͤ����Z���3p[T$Ԓ�9o�%]��r5Wf�T����� �	�믽=-Is�W쒸q��@U��t_��������z
��v�}��]���p�I��P�q�M��,j�o��e�"�9�1!q,�\_���z{���[Z�� ��EM�2FD�<Ч����W�T��2��jH6�i��:zTg#Ðlw��j��?���z�!Rb�yu˺�Õ{%�"(f��d���v{H�.U�` wˤ4B��'�<)a�)'��4CY����Y��WAQ�'��΁ߠ�C�h�5dS���w_i��;��y��EN�/�zH�'��H�P��vg��j�(��-��+!��p��	�ZY�/�<��`)O6@G�_@$��e�yHП����N���zpM�#v�'<���v>g�'����������۷r����mV�� a����߯����
"���_Ӊ�zǋ��:
֘\�B�����J��U��>��x�L���0"�0��X�9y��3pf&C���v�$El�	>��p��]�)�N[�J��D�B��l.��*˰0
!�i55t�����Z��V��[ݹ#fS�I�5��b c���������z疥Q�I�ԛ��>Ǉ���Ҫc��P5��E���f��R����r�a�����M'X���q?H 7��6.����V#H��:FD�R���e8��]������kb2�򅗧�{[�8n�&���pX~�����$@�W�M|�ʽ�I��ir!��dCX��.D�%���o.�ov*�M0��e$R��^��0��=��t9��!B��3�[ӈO�hrN+`��R8�����Rc?���U] Ti[�w���x'��h��[�i���[��Q�#��5�L�Ι�hФ�k՚`�R^�8BKP�^���+�q��s3`*��lJջy���͔:#]D/���ŵ��W����b�y� �')�q�"��eNkhX�A��l@�6��u��\�8�A�wM�����KZCI!B�ִ�
�Y%�=�H���H�z������|�-<���&*�I�!�+QaS'¼���Bf�j�^~XA;{�Ӆ����\P�����vNJڭ�����?�ѵl�c�ʐ$k)-��g���۬�*�ʁ/�ɘ��nN�W4��}"�nܩ��Cmv��)�=P�:Ϗ����p
�X��
����W��Hi���nt�>톧�iФZ!27/���[}f��������.7:��nt����K����#���B�7�b�����c[d
z>��#�'bF�� �\G����@нի�4��`*ax����p� ��R���q?� �v���j&]),��u���c8q��xt��N��r��SR�AU�V2����kޅ� `*m){9������?���#V# ��/Sh�sg����}���.
���2�x���Gݞb�B�O��9G�|>AHZ:s�lW������n�\_4��v]E�󁕘�*�+��)	ֲ��Kn����3���\L��b�7E�b��G����:̿���A��vbhtT�:��'<`���R�0�!Ňz�i0��Z�D�cǣ��"����h#�SYo����a��t�\o��$Y
@��ۿmڎ�QO9������D9a?V��	��^ЧXm��"	����}aXe;O��b�,��x�t�T+���">�-{�~�W�+��w���z^�¹Xꡍ}�|�c��p�1��C����r����A�M����,�A]�
�?n6�X �|�
��gKa��m��&�?�v]�y�:���5�i�Z.�ùծ�ͥb�o����A$-V&I�_�9�֠�e5�=��a T��,վ^�ii�g2oJċ�S�k���y/� �u��6c�y�3�y�xz����һ�@��=`ޤ���[�V2*:f�2�֏C�o���A�i,e?�<�I޻�a4��k��|1���N���ax=#�<];hE��R0����ښf��q�f�]�n)��T����g��`G���v�Јu��>���ң_V9����Bw,\e���X��w���KI�/o�V��m��@{��� ��sTZ�x���UC�`өm8u�
E;����5��e�Ů�3��2��k~��U����(���%@`}H���u�`�羽�Y��?Zv�S�'vKx�E���׍!����F��x)�tE4��,[c�� �y���^q�]F��s�·��>w�� >���\ԏs�B�yc*Z���N �3�8����[�ˋ M���
nG@>Ěa*w��c{IB�Wd�{I�W�r�����]����~�A�q��~\����c�0q�]HUp�,6&t2�1����8�Ǩ����,�fr ⮷(��g���,[r��׈�~?��$;b�I�����٧tN��y�ao\�w�^o(�QM�|A�|o�f�ۼ�����oKX�l2��1r�
)��_H� |��R�е�N{vƪ����!*0vz�����s�虞���V��t@��kN�RHd��*X��z��3%���l�Ҍ�˓LQ�1���0s�� /)Jo��v��ڲΓ;��9Ι(r؉�
��� �����,v��Y�ع�Ajw6����w��}�������.F��+���%ց�Z��)7G�����!�W�3����J�����k���r�P W�+:���XE��34%��*(1�ߪ/���Nw�� ��QC4�R��.A�)9��& �8垭02!"	Q
�ʼ����"�KM�2iɘx��6J�ѽ�3O�A��rF�Y:�R3P
s�A<�ؾ�9k�|�{D��)i)��/x���5ߥ�X�R��07�G���Fx��k�`S8ކ��QH��*�&��W�a8w�`=/�$R�')�����S4����\��	6���Z�X�dl�b�=��*МJ��Ÿ���)��=������D	�D�<���#�'"��S��G�P��&pe_[�� �F{qRm�u��M"�uպ�Py��Q���t���W�d���-U��#�A|\�
f�t�I�L���Ea��"*�Wd�[/aG����.-��mđt[��ܮaQ���y���8�
�hv�Z���h����&�wE��hHTo�]��cs �Q���hBI���ڼ�nU�2�Q�嶁٧�"0[�_�ǁ��^��3��Gg��gۖ����]�y l ���T�A�eH��x�eg�,�+�}�[%�HQO�mO��)~V��r!e�ª�M���T����g�4{e��%��`=�Ws۴�~VJ��n�S�a�ltٰ�'w�4;2��p���a�r?���;Գrb�����6T�����K����8G�2��m$A
�xP#���і�;�\ORfI7��~��{��@a��ZBڱ
9���W����균�����Kz�Z��E3cM��?�Dy��]�@��4
�>������Zmv(KǮ$m�!�`�#lČ��:�IT�/B�gDȌX�J	��#��P�pOi_C���m�K2a���"�������TP���O������Y��@I�e��?�:nH�/�}���x))-��c��=��v��@�W�A��Aإ�a�&'�!Ԃ:R���8�\�Ek�. G"�5���w(�O�Zv\Z�~޲�QxӸx����*�m�ҳ�3">qO�	�ir�2�����AAZ���ӓ4�ɩ	�8�G���%�⁷���θ��$ͦ`у%�K&?�G���ž�1'1��A��� $�`������7`×�$��ּ�03�f���O0>�y��L~F%Mx=�L�c��m����@K!�E��(Z�l�ic�^� �R�7�g���nQ�h�P�F��y��F��-<m:�5b�nV�ϐU�鐛c�yOB���'�QY�5����8�_�߱-�oֶ<�+�+�6�X����� �f�Mڊ��x:ɞ&]�М ��c��Д�\"�c�%>;��é�28x�ԡ�n#���d�cyϩ�i���4���b���g:u�����H[����t�Vݬ�*��:�M�[������䮃��I��Ff�'�Tєr�I�T	dz�H���i��V�Y(]��%r"����}�6o�&���4Hg̩��+�r���[ ��ǭ_��g���I��ay�f�7�-�F+=��K��@=x?P�š�փ-�LL'�=r�F�Hȷc�LJ(���e0E���:ӸF+	9N�K ��E&h[e@��]��M�-V�S�-�H�4L�B��.�PMV�fގ��-E�>w��A�M(
��aނ�V���#�V��'�n�s؋��o�\���r�����͟�F1�-],���2�͙����8;x�8J^j�n ����+��d�Bޛ��P���`]��V���G�$cŸ�}��o�ꘜu�������f�P�q���'6�?,��^� ��$�1�Y���'�%�e.xȸ8���s�O��l�e�&g8��T��+�ؿj�}�c �p4�A) �'oQ�a��8�y��2(r�w�������Ͽ>o�@	gY�Xs�O��$��|r!�����	�D%v���lf]�L��#�I~N(%]��s}��6���u�ӹ�s�3�c fւǹ�����K2U�K$0���	l�)����7Y���o�������sy $l�6rWO��8���>̄�h�uͦ8�S��L>X4R��;Ka�p		ӹ�9�/����.�31i�Ø�L.X*8}�:�[�$���[ݦ.����?��|=��XΛ}�]���= ��h�Ӥ�ˣR���;z�v�G�.�Qʨ~��)�?�����>���Z� �x.���"��B��T�8ڨ�8�B��>�����w�[b�*��G^W�~a���0����1�xS=6#��p���c�M$��c��kq�e�̥HP&EG�"D ��X��%��s�|"�7��J$��)
)�i�^�{�eH���M��p���n�cw�y�^%(��Pg�El��q��_跭S��vBڌ�n�;�3n��-��8��L���v9r/(_40�EJ�/�)��a�j�-���6�o ���L�ɯt\Ӫۅw�59��t7����!7�_�t<=s.��-���4�}�(���7�9�Ξۡ"��WT�����v�/]�R���q�����>��W��u�j	�@?��k�ȷJMX�/���:�����$X�P	1�	��?h=6W���RuWa*q�?�?R��n���Ķ��y7���ƫ�P:[��q��'�S`>��BQ��,a���N"�]�=�ՌZ�GBx��xU�0,G�����G��[h�Ž�id���3|oQ*�jx�v���f����<N�,��8
�=`�a0�ξ��/e���� Z��*b�����DS�io��=�Z�G:4��Y��P��q:���#v�5K�$��Y��Y��7�8`�:*�*/�ډ`2>U^������;y��i;�E�!.`�M���7heih�$�E�
��5p�b�n�\��-�;Q���ypy%��c�m��(�s��J�S5�ی�j��z�BW�˳�/�p�.����mp2���*;��qL�H��#�F%Axv3]���y���o>A���~$���=�����w����p}!�V��#?ɉ���ZXm��Q�o�+�cB���n~�%��J�?�|�l�]����]۞+$�� {:��}�S�#خe+nҋW��M�W���.q}�Cz6���y�����&Q9�=�(�Q�j��	t���>�8�i^�?b��o��U%53"f�'���k���-�H%��BAZtEʧ]��bֵ[�Ǽl���B�I|HhL�K̓� ��9��S갆{.��$!ë�\���bK����.C���%�w���?d��m>d�]���s�r�Z�sh����������� mD�W�U�/�Ψэ�P��W�I�d�)�<0�9&,s�
ZQ� �g�oG��P� A� ����Af��-���ۺ�����z�g�z�F�`9	���tx��7��bah`Aؠ���N�^ߘ��xx�b�7=�hiy�1���<w؟�7��wTuǢ�/Ƈul�8���4��؄6Q ��G}��{4�ehpDH'�(�H���@�Wrբ@~@�2��R^pw�F��Vǀ��e��
�s]�U/�M�L�18Q����u��y����&[U~+��xw��B>�����و�����'}�QD3��9tY9���� G�V�8�ej�O��fɇ:5;Q���Ռ��<�w�G����Z:05^�X}��t'O8������i�l�̌!#~"Rݱ���j^l������h*�!�='p�2Q}�H�(�"�(֞�����R�	�l||^�1,�vS�����3���±�oE�e<�ݡV��˖�#e���� �����9F*R
l�C2-�SqJG?���fK)\��崛F��BJ5�!�q�LS�Em�ed���4U�W�4"��]ذSC�@r����u�C�~����㆜mٺZ����00�~�(˴���!X~K)����E|(�e�u1���������.| V~��L5����ێ�@w����eum���K-�Bv��|\�ߛ�}i����g~}ZX�B�����r��=����Si.�����"��-]�_vQ|���M�+\��e�S��u[(��/���wA\�n�nCԻӤ`8���և���o����'��SA@�3�0`-Q�7?�[U�U��4���
���³�!�/:����Yh"x}�;��1!�� ���w]�vן��5A�#�oc���tNc�K����-}���)�9����@-�Ǖ�$}OuĹ��)0�.)1~�[eB# <cp���w�� ���1�P���4ǈ�Y��F���@�:3e�r5m���<�ul��sX�q.�;,P�Ԍ�~-T�A;r]��6!�eѐ����#��%>Ӌ���(�H��,�ŏH������:k֜��F��6�2���u�yr7�~ �O���[	�gZ��H�e����s��Hɝ<l���vf���L(��q��-��ѱ��� �]��w�u�L�*x�U&�6�p9ŊW��1?�5=�)�	b�0���C�b��B�5�4�27��5΄�'�d��3	a��d��Y�ϋ˷ ����=Vnr���~��I��9<0~�G��� ��C��-I-1'�4�+�.��yqJr���q��W�m�MD�0�41�DΡNh7��EC�MC��B6u	�g��Kw�K&�����Ob������N���ʷYp��e��v����;��&#m��=l����2�<&H)L

W`Z&��r��<L�1Z�͝����y�a'5�K"�/i+���)3��V�c�6���k���Egb�/`N�ߗ��'��ɻ��Z.��Fu2�C_R"�X́ ����l�rSJ�ͱ��ê�S��%�i�)n�:�-�ɚ� o :G=�k���<"�!_���N��ߵ-^e����e�$��VAH���c��#� T�'}�����˟��!bR�>�-]��M��KQN�C�I���E�K��o�y���i�j�l�U���R�}�NWJ�C�Y�7ù�1֜��"�G�Ep=����JHT��W���׍�����e!� Amq�j�^�X���:p�̪�l�����QCH#�m�A���F�1�\�C�Tu�8����^�<N"�b���DG����0x�N�2єB5E�{�\kc��K:���4�P���˝V�Ҧ����v	ۛWْhY�LA���v����i���ۇ|H��I�3��E��ilJsC!�&��SO͙/�"���*���qs �8w��������i�k�7�C@�mf��Q������?v]�����O���U�Q�UX�9@!��� &pm#:�'�_`�(+�e�\��C�F����6c�1��gӥ9��Z�$&�8(������m�g�ݫ+�mK����� mV]�]g�9�%_N��/<'&Ŋ��2g�ZUX���&�h�}�,��`��2k��n�	��~	:aRM�sS�m_I|iQ�����"朋���A��7a��@�bn��p�pc������	?�.��Y�f��+5;HE�%,?�x�F�$X�jlt::o�$�)��I���1ڀZ��K�:#��[~��X�W���:F-:ǚ�R���(�]L�U����K%�㘝��̍���o	����v>%f~���|�y]�Ey�:�t����S���.}�n7�G��x�LfnY�}����n᮶k�M�M�	S�a��۟;����L��)�L�	Ȅ�#1~m����u��f%���K1(#����Ҹ죃[��C���m�g�,Yy��!k�nٞ�CBo����_�L�@"�U��k&�$�{T.>��oLa�j��:r@<(����d�D�Y�)��Q6� ��l���+!Z�t�#vږH�5(���vҢ�0��
�$��3�|\��e`���qf����j�.��)�~�lۼZ����z�wWÜMq���t�Ixd�D/�&�����o�N�J�z��"*�QC�H�h�E�ˍR#�����G4�X���͛��W��W����	ϲ�$*��q|B���E�.	��¶QÛ�f�F`�T9}�>,4d3 ��|_/�/�'HK�8eR�a�䣙f�)D#�K�>�p M¯E
�nuf�����o�}I�K��f�ɉ�f���Z.����	�o�$_���o"�����ad����NZv�5ټ�;��J�߶����b�i�H�^Q����Z�c�	xRP���׋��!�^����b����'��'#o����^��'(0�=NV$��S73+?�u��j��n�E�|sf���K�hw�am�0�x"����d��@4����(u1�E[�`H���,*�G�b뇬�1x5Pп�U_/��ͬ)���
������ud*��3���Ŝ7]�1�v	J.h�B�{�#?�=�X���al͠>��D��6&����Z5�L��T��W��a�ROp>�, ���[
�p����o���c~.L������!Ag�����+IU�(p�v&��.�LU�#T�N&��S��f5VCJ����R?��d����"��)�	���o�>_�n�7��%��u�u4��k�Gb�M�
 XO�G1Og	~�)S��B7Ot�k�s��Si۰Ϻko��asZ�mGPqUՁ���0��V���w� `��;�O�Y@�ST���[�����<ҦF�6�땔k�z��C-���Ih���T�i�[PSɀv��l �LYQy��T_�~\b�IV����bcX��٣e�b]m�iw-7�#�Ws#��L:�(Q��W=��n�8��_}��c�-<�M�!f�:�U�\"���A&�>���C���X�_�GT��Hg!�~Q3Avr��)]�^3v��޷�U/���U�+�e�lz������2��,��|N�R4Q��" ��X�MXM�\�X��C��ɧo� ��f��iv�{e����y�fI��z/����������5BI�w����U�w��p>4=қ̀���x'9��Lb	k:b�,�m��'n����fD[����Ϥ�{��`�{+G��h��j��W Vh�7�a�-��:3����Cv�{]�븍�Mo�W��`x
��˖��Y��M� )��n�<�o,�\�e�y�	>� �(�Z]�=պg�w���=�ް�N���2_�f�^���=�SY��N���Cj�̇��>t�)�P�d�/�l���L^�k
��6�Pg���tg
r����m���J7\2�_������2��{��/�cU��nﻉfڥ*��b�L ub�����zՠ� !-�N�3��64������.i��ʌ6��ִ�&z��B�r,w�ؙ���^~Leg�ͥ.́��M#gH	�.�j�����b-�;��'9�~��W�`�g���-�5�f=�:.σBc���ܮ�j!�S�*�C�\���( ���3yP��T�����T�c״ߑ,!ߞ��J��Dt���!����gb�~)RD��_bb�5��)+R!���NB�F�n))�,a����\�⹪�n6$�����[#�����y	̧��e0ܛz�$�x�<w9�FΦe����*
��[�N�!��Dֵ	V�){1(EMd
E�X�l!�����у��Z;��g3��[i�-.�m�7�+�j�&1�?W���Z]�<6��s�03��V��9.�cu�U]��1�\P
�����rģ��f��v,�=X�h[}NKΨ	�7�o��R��NM���'�>Q}-k
��i��U�k)gw0�H��|O�b-����C/��p�~�^0���Tp��v�Z^S-�+�z�6{��pF�HT��
��2iTlMu<||5�b�����BS��g5�����Ir��i�4V9���(^���b˱�>@���j$|����. G��0��ʣ#&��R�@�Mv�a+������揁�JO��_��i#��1
���p�4�H��:	�P�E�r�Q�jϵ}�醖.Қ2�b�����S��O��m�dƱ�X��SוW�	�0l�q���nU��K=��Y��)������ݪ��(Ci�s�ߤNo������;/��\yr�<"P$j8���W'δE��V�u����6S�;�̸.�0�R���=�py���F�A=�K�8��Oi�����9��"z�~����L�A�E����	��0ݪ�w隼_�I��q�q�N�5O�0m�Uљ��R��������"�1�6)�X���G;�Z�b�����p���z�=�~"�:��`	icM�R
I�b�%#�p�b�� ·er�˘���g���� �>�2���f7Z�J&\�r�Kz����-�����j��n`OC�uL�a�P�*�i��:�lH����{M�����i@�1R[B�s[93W��P}d��-�ȝ�fn�-�Qq����\�FW]�5m�&�޳�(��x�BP|cb�h�o}��k"��7�Ī�����Y��#��q���+�$�"e�+jR��|SR���)1md��jN���˝?�UR� $w��N�R��ij�N�?�Ɛ	����Ÿ����lA[O��	.)o�<�y�bb�=��A���n>�� ���a�1�UX@L��he�eTa����)�S�X%w�cj�m{<5^qP.���|uӪs�C\�	��T��Bk33��^�n��J�k��\[���G�:�����d����Υ�s]�$V� 7�Y����ZS�+ʾ���1<$��9_��ݴ[��������k����G V�H=s�a�u١���(?�0���W���[�}�o$kzd�ਤDk�F'��nW�_d�22�ׇ�wX���n/�w��u>*�#�� V�6�+sԄd�����▵�R����65��C�a�H✶&G�A�$�qI��j��8��aWzf���gZ�q!�(�uX�V���s��T6���&T��zk��8� A�C	$��������תڧ���1�%�{�y����x���TQ�3䌧rt(�%�d�4%��|+D8Zb5F!����(Р	����9 M'v+�|�@��s���e)Mmj�P�c %����jEf����g�vэ�3��
�4� �����YjS7������``�$���F���i�8S�e�R��:(��".��}�G�۝R�˰_]V�A��U'��"���'Vd^��لE�\\����ܭ�]ġzݓH-�O0�
X+DSS��Вk1�ʄ����K��)��I���Gq}��
����x�y���TaJjOhW[��-���S�8d*͙����{��j\d蓙�U�n�󖌦�P͖J�y)�Tf�/�˭�<Ĵm��*�?|�p�"�I^虐���yO�{����'E+M��� {Ϭʤ�,�H���R��>�P� 1��l�e&�L�?�\�V{dN�+���4�	�d��NADu� ���|�ǂ=�f�2��"I]n UuVe��i\��8�=�����<���RY���j��s�mxWB5�_��X�20 9�q˸�p\�_i��ލ��K�r~x=���*A	�n3�U[�@���P�YJVw,��7K=w3Tq��iAeiy�'_�:���Р��,��V�p3��k$!�vH���gB�i��ɂ�)?�����Rb��<j�L���H>Z\+�2=��u��z	�ӛh݅8)K!��5�T�xg��ƽ�S�m�/Z@֠[�4̰ZA�Z�:_��<������t`�l�?V_����H�Hm���$RF��m$CYR]~�W*H�8��"7IU��W;AT#�V[E_?�������'L��tW*q+��O����h=����v���:�Xpc�p�6$�&T���[35O��C&H���	�Xf��Y�}��kX��J�S��F��PJ<`G���U|�h7P��׉D��S���Ht
��Y
j��	�\eAdH��}����C�mYnʧ����q`�V���+l�O}\�3��E�I\��0C8r6L�|��4P�ެ���ƭ�)q�x��Â�8Ҥn��ѡ;z6�ua- ~�jj�P�W�	��UJU/'�;��� 50ڗ�QEd7�`�?����ARZ1Q��/��=��@������kAk�`ܠA6*���-���M��8n��V�?��D�S�>��VZ�T��`��!#����?ͳ�(~yN�Xx��e=�ɝ���i���G��s`�;��p�0���G��[G|�����x'Z��b��x������I����}�MTFs!	��k��2��K��5aDSIDB��&��\)W�IA{��lЇ`���܅>2j����K�ًU?��8�DW/2|���AH�)>�[}A��V�4�6��6e*�J��GM�k�����|��`D8����<-֍O\�" �f�:��\b�l:��9��$�#���{��S%/�������J27 �md&�p������Z��i=<����c<V��	�ΪH'��!��ui&�6��m��wbo�ySQI��dMD���|^��X�>RwC��|ER�
�����t�(��.����u�[_l�m��p�"x�����'U`u�������¸�w����)}Y�UӇiO7Q�uw��������Qj�`�W���(�\�>���x���<�!,������ \v'�D&��ݠL;�*_lx��7rq�\��f����)OOoC6^�E��T@R]9��}� �¤tvZ�uܟqτZU����Q?��b�U�`�ԗ' C+y��ω��s��Hj_�&�e��vEv=Ƌ�m����d����(�y�Z12~�èC$(���e{ΗCmqo�O��H�9E�D�
���辘9�+%��������0�:�p�'J�5���V��>���G�.^E<=��m�@.[ϒ�#,qr�T�N��G�n���E�¬�=���
|w�s���ln:`�{GUꛩι ��q�WVvq�&�C���J
>}��L���;jM���{):m����{� D�+�؍�w���D.C@A��*��Έ���^�9�dc������!P|�՜t���.Lހ��|�:i�;����}F��m����LL��Zr�,���^���!T��F�W���/��[��V�!�p��������e&eq��d���]~<��X���JSp#����G6�)zv����n+��>*���i]/�֞	��q���g�t�n�\{dG�xtX�z篣&ֈw�0����W:���؊�Ǝ�75/=����q	��rf7���� ��,Mk�M%10!#T���-V$m�(Iv�K6v9k�)Azr$'�v7� �����K;�5%:9��|��<b�\�ଳ:� ���j��5��l��p�F%d8��0z���S���ҡ92�Ww��O��or's�So7�?|�`C�a�΋��M�/�^�t�!J������b^�	P(�?�d�<"�E�o�]ʍ�{�y]��]:-��6��p����7?��]��Y
.Lv����]����Q�%t,�ư�h��C�#��`�%��7ܠͥ锢+֮j��u��u�.5�`��g�����=�����Yp1�0�?0�W�71j�tX � <I��-�i���SV�����>6���|�Μ�\����dlI����)��IH������b�Vnk���(ҾS��q�UB����S�
g܅ݹ�G���0%C<ge�4�_ɹ��U
d��Ej�l����.g�ZK}U���}�z�%�{0#$��zt�VE��(���E���ɍP�(�?R��.1��`��upU���;'�Î�U�"@e����[�8��T�����nvw��Z8[mtĖ!��5}��W����bM��yU�e@��Q�"oH k�?�:�^��k�*F��>KR�M���_s�����[��фi��q��ym�:���BΣ�ʧ�!�V;�J�Nם��D�9<��de��5�wZ��S2�j�m�ۦ��0��;��l��-�r9}ՙ�O �bhY��em�Fď.�|�`B��v3^"!�VE�TN;�����
w�m� o}���{H�I�lȀM�|9�j��������~b�޸g;qz�;{|i"�Tulu@�����j��̡������':,���a�\e$׃�JW/��Y�<�Q��76�A�u}�W��'�K�����9�)�]Q��
��r���t��ʝ�埨m�M�2���X�%ߗ�_��x4%��o�\7(�u�	1�� f7W�����yK$2�	��lh�(#�+�A�Iɓ�MUUKJTR'&_0�a��#�{{�{H2G[si�"�,��͌op�3�b:lf҉5,l�r��v�t�G��i�ꁫJ���D_H��V�X�X�^E�z�A��M'�q>1P�LX�(%w�DE�4����9q���(�4���J�C�q�5�vlC�x�&t��;�+H}w���&<��f���JY�f�wf�ٶ�/�XH<�rv �z�m�A��n
'vGLd	�s�Q�>��?��l�fn�W0�jo�Ngޕ����R�	����2Yjֲ]~�q�ŕ`�R
<�օ$hS3� ��$<��po��[��W��#U}XzM�_�i8�����u0S-x�Ek�CgIͼM�� ����1���Ӷ>�:q�y�����e,�6 -j������(lf�NKmި�?��ҟp�S��٪�8���!�BY�$*,V,��2D���5����bt�؇�icF6�M
|] C�adw`�Y����6�&y�����t7(�|)��h	x��?�t(#�`~�*��<ŜB�o�S����*�)
faz��Z�{��}T�n�Gb���z�.������Ok��A�*�D����e���2�=,"ox��H����1�e@ݤ�s8O8E�������t��q?11�p6�0�[��U��7��3�N\e/¦0���g��&.���>̊������ac�^�����!��Y$^����S�%��݅jp(ԻxK�����g����m�q���-�y�z��j����57�����;��4:7�N����ҦP���+�'���.(+@N��5�򳍲��|�ך����~A�ƕ�~]h��J$��S�'��n��r���5��W�-ѐ1��2C��eEx^�]�]�]��.��y���z)C�A3������&�2�E?�z�ޔ��o���:������O!���:���z�~�w���6�v��}�����F�tg��T��*��,���f�)O��x~AR~)wG����Z��?w�E�2��o
��s�3��x/��1sxH�7�C����0����_Ԩ�m��2ѥ�qDj���Ԁ��})���[Da�t�g��DQ���l?)�X�Z�7�j��81}U���%-f[��o��q��e�a��ɺ����D��H�K�hF�jj��Q�%+����	���*A$��ݭ(|.��%���}"J�+����~G�ÿ]�X�z�80�����N"�6c�6���x���G�]��P�s��#n�δ���M��v/ɲt\�-{�O��c6�(���@��d��Q[5e<��pwe������cL><������b���
�7u�P:�>�������#cY#��+�O~a��Ѹ����e;'���}�l2��ڳ;�Dp-����<F)��o�`���.��H�(S7�t`3J��+b�)�F��>j�p����2�S��!��Б>��bgA��;V�P�>^���k�=V����t�G}�al��N��ԀU����Ńn��Z�fBO�]55�_*�Y-[��|/\��^��ؕ�#�z�`���p8j��}X��4�����TyR]���X��I��d������c��b˺�	H,��S�5l��d��w��KlQÙ����uz�]��]��#��9G���5���)��U��RB��:�z���������)��,�7�°b�r:P������OD��jc�B�-F�@}�ӷ�9ގW��EZ���)����ޕ���]R'�h����m�%f� ��ޢ@���E���I�;.l�c-���AL��!�ef'5�A���<�Vc���i>_��z�M��L9��%�1�~�s�p��0IN�sgM/P��`+Pg����P�L���H����e�!�<��ޛ����RR����9�uo�s�����N喞6���E�����1MtaRc�'V�N%dg���7�YuT��|�m�:tt[_�Q_�_�ƚ��&=@r��!ݝ��kю����?��}�LG>��I�(S����ԨZ�{�t��cbz�����C"��z7~ʉ�W�l]���]�ǒ�����1������{tlcE0؀���	��^^������h�V��*�6
f��wC����>#����؝���Ѕq�OY������%<c�.XFr;�FC�E�hP�	bUџMV�!t�}��+�(�<uh%���I�9z�;AE-�k�g�b!O����zR�ÃY���W]��Z��/O�(G��)�b�ǘi�t<�Z�耍�O����A"��!� ��\�r��mk�qS�8f�� �0 k����A'��AZbO&ƛ����w�G�=x�8�d�l':�����D�h�&�����~t�mij<�X�R��|�Ue	���q��p�M���i��u�� o�Lr��|���~�S��/ڼ�@�M-��4���sC¢t�U-����H�&,P�Kg�;��� ��֣�V��&V	�@��L>�)��t?����P ��վ^��-���dE��W�A�!��J�}��"B�$A�)��ڮkq\�U�0WF2n_X�=*�^���x�{����J�'�O��R��42�Kk#�-D���_�N��Fq��E�p�Ut�h)y.�o���#��?>h_^�������`�B�b�`�,��)�QzF9��z�1E�/�dN��_���# ��%��-��Fly�׬R�����Au��2�,fC7zU�݅T�J$0)r�/j�X�&3)�ŹZ�D��9�L1{:�$�$	1~�:Q� ���jW
�5�;p����pg���v�B 8ң������ޭf�N�[��0�^N��?�)Q�f��iI�z��%��u�7U�����|���AA����a�������o����{�uYOF��|�K9�C�xdr��L���Nf.�Ю����_< ������zz�|_0BI�$7�:�WCt�PA��Wo+��Ցg�\���A�f��>��£.: ����t��;�f�ԮK�9G�h �Ϗ�&7�t(%T��c���B	g��-w������J�E�=pr����Ԯ���N�|3�I�K�۶�CAI�۳BAK�Ci�4[��,o��p|�$^Yd�ע�ЧS�` ��T*=JHU�g/譵TBi��#��s?r9ը��ESK�%�W�۲Q��M�������m�h��9^Q��t[_�����ďM�����>t��q~D|@œ�F�9�-���g,+^��-��H��Y����}�@�e�OX��S���nAA��D���Gs��M���Q��д�'��\�^h�5�P��?Al�a�z� Ĥ%a<���'.�8��!�%ׯ�1�������^ʛ��6'$Ev���Ɔ�`�=��/{�L(ļk�z�tPt�j(*d�y����3��nߕ�+ݯHFLyG�=�k���|��K9����t]�fo�c~ ��XT,?G׋�i����f6�8�kc�a�L�F�*)U�B�ܛ�eM9�yt���0\�:I�u�L�o2� ב�ڍ�C<FK��!�4^Pd"E�r:��L��a��3�R)��X�/��< i���~=��$��)�10��m����s��!�oR^�F�L���Oզ/ C�1Em�-����]]���J�n +/>�9P^2D�g��0���ࢡM*'�/(D�;�n�/P*"D/H�ޙ�"s_�Z�<$?*���n2Y�=�)wC��Su�b�i J��LwN�wO���}d�vÕy�㈧�-J�<4ۋ���W&���E�'f����	���6��b7��;Ju�+���j�Lq�CN�RW�菇D��<�ZI.ذ�XA?�4�!R���8��ZW�i��0=�Uu�ݍ�cƻ�2���0�a�GM �M�/�0:H<n[����A��
.��
�r�����W�+`'T�H����L��A�*L�Fs~���ǋ��tH(]e��������mYЃ�]䱽�EG�wKE�K��r)AL3���~�h{\S=Y�ۜtz��m�Qs}�8o,�1���=��¼���p8�=��z=�ݩq�62�V�ޚڼ��ӡ\���A�Hq�i/�����n]P����C���d��%^��&n�[�М�4�����������htKD��n�C���Y���,���i#jL��/���I@	1��ik��2����xey�T�����
F����'и�R,H���a8�2�?��V�߳�1�_��'X\�*���V�a@�e��u3����P���#��$�C����!+�B��P�5.I�D��HD]Y���p���^�6�آ,���ir���
�׉+P�eV�W�Q!:�NG3c"Ⱥd�"���h�<���%ǳh`�x{�g+��8hz������@7�h!Q㺐eS��OÕg,��AZb���wH�S��Q��0��G�Ma$
x��g��8A�1�5���OX����C�qT�5�(ǒ���E�/x�F�p����,�����=�M�  @@�o�ˬ���h�XY:6����a��A���_VV�"pȶ0��"I圿�zX9��Kl_�W&�X�D�r����/�S�o���B�&�>���s�����<��T�K�R�.��pm_3��Δ/,��HC���_:M��?E�+������)�z'�rz�_�2�'�����̎+����4�?��;3 ~����>�. ��,��tR(�e5�� :RSxk��&�@��2����e���bE�F 1m���$�V3�b�O�H���G�:�	�UO��⣀BU�܊4������C�o�w�ʖ.|M��|�x\�,b�^F�15�����_<B�wg/�<	ӝΫ9�4�Ȋ��~��N����F���砬M
�F�Q�O�� ;�hX^��l��h��I��$���7�?���)�B323Yl��55snҁf8[=$@�*B��z49��h��]G�Ԍ��Y��ڜx�],�,1f�]��{n6�#����?q?gj�#�28��x��N�f�72 �p<c=�4d�d�=�ngͤ�H�g�by5��'C��&�u9D����ذ| �D���������@ٴ�O�KmR���g��(?txq ���]��!?���>/��
]j�?Z{�xT͆<���0�S�1ږ&Z�������?����M��t�X�A�c�<�����/�%>����������"ȯ��R3D~�J�=� +�,���_m�۠wֿ#�\� ���.5�d^q�E�2I��L';xR__ �s����+�O;a��AX��E�����0��ĉAd1�q@���^��\7]<�|���z�T��6z�k��Jj��̭F�-DZ�S�0J�b6�m��d�"m4)i�y���4�?fdn��ɵ�	�,
ܨ�0����6�����Ȱ��Lj י�v��D��-t���A�aHx����]���;����Pb�s=U�N� 6��Jx%�Jv �e������%�D��Ddb��ɥ������lI�'�>V2-W������9ad)��V�iOS��&z8D:�b�ھ��W*)װ'�^h=��T}��(�,ΏW̳�蚝n/F����8M�V�^uӮ�7t���6�b�u�6��AO��Q$��٫��A���Ų��n�K ��a�o�]hR�U���i�5�J֖q7����R�"M#��cn��E}<�ʉ�	�KDu���8�&Ů0i~:o	�r����,�a��y	��nL>|�UDa�N��ޯ���|6����.����Զл��*$��뇃I�"�����[��V(RqK��C��m�劆�=V@<��p�X-g��`�rC���Wp���Zɇ�b�ǯ��F;���%g�C*S����ק�|��s��oz�h6ZL��{~4^H�rd��"�d���_[Ύ������*8:vwU�˩cv"0��d�d�~�]mGc�V� :|�0��r��va:�!%�����{+�Ԫ��с�C����˫��u�C잳T0^�~מ�F~�vH�P�Y�/\јu��I�BWm�- ���'�LI������T��#�P�O���磘Gi���v��'TL#�]�R��Q�
wV�D�O��W���͡�;���w���+�d�fs�&>���8�R�Ph6�$����K�_Y�;�M�ED9����lnlA&��>�o,p�X�%���3�1I~ɷUm�,�߃�>}������/��/D)�����=y`E
d�uAʱ�W��#��?�'�G���s�h{:m��J���[﹅�I��:�������*a���XÅa��Ӊ�gѩW�+5�דL�G��Y6�h��c�T�͑�q��N/��?��gD8a+ha�*���{��!��r?y�iq�����x'��hq��PwU��}���%�����ƚa#j�����b��WN��ߥ|9i/�����=�p��_�lLw�^9k�E[
r0��Xd,[F�_k��{*���vզ�m�qEl���~�I�Z�H�BK���o���H��cn��E*�2 Ү=�U��:�l���т5����bWyl	,�JTmj�z�3�Ad.�oq��s�i$S �(SlNg�NZ;EJ�����:��IK���(�a�I����
�aM��.`�g�8�IT�Jŕ��K|�g����C�qT�RFEM��Vwl k�L,Q��d@W�,S�n@��J	���DO� �&�T�+�y�/���1Qk����㑐l�f�Č#5���c�`¨����h���8icFe7|�R������A�Ғt�H`�����s���{۠��$7���0p�ٿ� }�&t����¹�fA5f�E0�V�Ⱥ!KHgAL��8F�@!80v�CG�j�]��'x~m�#�T�I�{�:J0�
�q��<��h\~�����"��Xz��1:���tg+Z�h?�)݌t��"*1���j��$A� D���Y��4��041�;���	=
���$��7bƾǣ����H!���(�*�u����^��:��a�ĳ���D^?�ڥ��� ��Z\
i�39~Z&�Rڈ�9�`�&�΄z����Ј�-��s~�[5���Q��L(1䌐,�5al�t�R��V�Ɏ������gڰ�`,,#��?��,��2�ӻ�&`�fY�iV�g�*�2��&��#%U�G����SW�I��""�n(�d|��>�Dw}w����G*��0.��w1a�x�����C=bzXGh>�>FMvP��.4K:���B����Y���gIwT�*;_R�{�	��!^�K�i�>�.i�8T_	�V�z��!50����ý�7&=^�Y[���hG���K��k|�k��{0=�EB+	��»&���'M��c�H��p�z��Ps\���q���9�םǟ0�6@X�]�0�������l�;��)��5{�`��zNF��0�v��trF\��uOw��3�UrH�Y���	⦃�_>�u T3��"�%��&b���
W ������5�Sz��d�&����?b�b�7.�G����U��B��dg;��y���.�d[�ج:��[w��B���M*
���e���DT��X�^���Dz;�#�Lþ��@�4�����ܹ������6�-F.�)���E�1�5��>]LJ`ԇ��J���nj�g�?T=�J=��BQ������R�>�Ɉ��meH:{L��'�AW������ ���*v����t�<Լ4R��x�z��|c�a0��j��a�{��V�HL&H��W5�����^������[!/�=*Q5!&�t��4��3�����K.[�Z�*X����Kӻ-T��8�bj�!ގ�ko���&�2�l�T)cD��8�!�����r�,�㖭������t��!��S=3il��YA<�=�/�X�o�봁�*���1�C�Sݩ�̩jg�i�Bs���l^*y�?�㮜e@���,�̫b	V�4�6Q�#z!��:�����ԍ,/��H�Q�ܧ�tJ3`8u�u�v�h葐���6S���{�x+� ESl�v�f)�V������(���D�b	ۻG$+g�q8��^��I�`y;��>�H�L.i�(��1KiJ��~aK�g��[[�&Ԓa��3>u!�]-Y��R���ׯ�:CE��l��O�]��H���Y44��=lp``ɺ�
����T�\����;��N���
Q�����4Z�$�΋]������s8x(rcd]��-��cS1X�kF8m�'�����
�y�e��3�����)�4��*᾿�5��KFb��9e�8�����̠z/��*~%���}�Ћ\����L��e���FcN�Ѽ�����zH�?2��.�0M��|�,v_I��LɅ�>����-ߧa�����
B{���B-R���os�����S'ɬ��0��Nq�I��&'��Cj46k�4t�ǻ�W7�piAcyu�����X�b��a~�� �c",<��ɀ���ZR��y�@}�	 �5��B�K�_@ѽ�S���p�0Mū�K�,�����C֢r����(ɸ�:\ 5�d�h�t(�zû�	nYb�C ㌪��^�����1��<���2:S�8@Q�H�0�NS�a��3���+���)c�G=��J�Ԫ^�n����J��ѓ-����ʘ��Xa�e�c����̕�+�ԁ�iQ�"G�#W$���0�[����B�b��[6{<�%�ꃹF3���/��j��q���u�7��g[FY�k�������0b9�y=g��۬�G���7n ��+ޝIB<�u�*`l�}�������d���b�5��_�/ ������ư���x�t�w�l8kpE���@,R�R��,�!]dU5ݤ�5DB���>����!�l��S���$?J�z��k �Y,9)TĻ�ٹ.��>hL���u� �ˎj8�������]�1#[H|ٺM�F�����搗?Ra���%�����KC�u�3�*k�-��rI&�Ey�PF)�G���MUTu ���� �-���|�+�����'���=R�@��p�*A5~<���� ��m����R|����q�D�ii��n���U�?*��0dp˂�+��E�t�}nTݛ�qLG� �p$t/�s7��7�P�T�ϱ(�-����j"eq��X�B�*�L����ܠ}��O��|/���;�Ҫoi"$/��j���j0�,�˰��"�������'9S�񒭠�Wg�DL��	)X�@�y;��i�N�I��S���m�c��yPh=���ao�X�5�2������Z�ϭ<�*�O���N,���[���0�Y]�I�lT����J�9��)gp�}��6l�3�+7-?�X���+u�!+���\o�B���lVV�w���\}G���+�h�6�S�g`��"��s��X	x��t�"2y��ZU�z��7FR4R��F�w����J�J�^#;[(Is2|5��n�2x��Kdt�'�n$�1�4�.�V)|�-O�mV��e�̕l��ŜGGV��GBu�ž�Z�QP��L����@Ŵ��j�q'%��&�@+��*v�2�%q����dl+����N����>pvv�	�~��.ѱ����%��R���6P�a0%[C�":N�W;�Pث.�M8�w�����?����Sz���i�rvڃ�#�Y#�^���gTы!h��8d(.�^�u�����r��r��v���̏��;0�'1�/j1�+�sZ���������1�����sq�>!_-uZg�D�2�fF 7���#�e�^>�_5���;�N�
$��eE~\��\y�0���I�C0>�֒9�2b%�{A\�����c�g��΍���x��?���)'v`-���c�2�u�WP{9���m	F}�8���.��,N��܋GwZ��S�gjl7�x���О��z�����(܅�I2����	8��V�Oa���!�0⑲R�V�8�48�+�_�����ʥJ� ?���*g��#(Y��Ȋ42o�:=1�����U�gwk;)w����U|xKMIs��G��X�V��7��:a�\��!0-����#�uyFQD)ߓ�0�Ų�K.�8`�k,�]V��QuO_�+#P��-�'�,꘶�R���{��O�܀
��� GD�I��Js����4��!�@�=x��Q,MU�2�Q�_)8o���a���6E����Jnvs@g��
>��>k�-]�):��i�7�ff�J��l@��b�X���nR��w�u�/���?&�}~�����4�K(�|a1�z���$E�2g�A~#�0�zdفL�Ƭ�T��w�����<�n# Fb�֘�੅�-L��Jx���G5��>�V/�'���#o�=���b��g���Ԇ�Ja�bq�����1c�Hq5�x�|���0*26�Q�$X]�z�E�|�Y:�����%>V�x���CL`]��_�p+1���
6�����א�f���ή�Q�st�X���5�IM�5�ڢ^�T�T�^7^L���8�]�$�Cز( z�4�8|���$\/���\Y��Դ&�8*{P����w(�$*XA�d����is[�Ԧ0��{��_�"�ӟ�3[�Έ%����2,9����\k�L�b�@v�k'#�)wy�k[2��p}�4M�(z�ok�vA�i�~�ȉ��x���-�;�ž�@���p2�F���sH��U���b���)kK��i�.Kt۳��ڏ3�R�*9/��𖕶�:p0=��ې��hc�E�\��oZ鴷��QD@�'�R���@ֵ=��N�I�K���cb���yPh1B��Y��^W@e�j�it��������,�{�dlf5���"F��I4�5����w)K�%���lLƱ�l�Z78�*��/�6Jv�$���U��Ë�H�;$�u֛�
��wJ�L$�6�˴$� �O�ufh�F#z�o�U��w#>G�E���UH�f�n�ܾ��B"�]+���eZ����MM�:�CR�Ϛz����)�u@i-(.�m�yv\����)tU��R�>pt.Ξ�N�z�#
�M�Ĥ���4���
�!bDwK�T@&~d�R!�n�ռ7��u�����0x�^X]��S8�̚�VI�8���鲔��=��aQ�� O4�gk��vEƥ ���`g	%O;�޽!�#�,o�z� ;��)�sx�ǁǾ���OQ����g��ܬ�n�\ l���������c�٩����}�ț+e� ��?�z%Э�T��tg��deG�|_0\�2zw��t�p 8���[����J� �/Q�:�AH	��w���%cp��r
���1]D�n�t���������a���)�)k��,,d'hO�F��m��}��q�}�l��[��MЇ�P�h,�J��d�!,wx' �Tp*��Qd��LP�z0B����K�(>���2Sq�ެC����!{(����*q���R� �Џ�o�^���Ly��K��j�B���,?������v �«t�
�s�h��<;��#���*4K� P�_�b��A�,W�2Ac,�*��^�KwU��N��i�N��o�/�q�+]�P�;W�����L��Q�8��^��H�s���\�vc��?^�"���`s��֝=T��e��F$��9z*�/X�k�O����P<)�L�,���f���uTG4�%��eSΣ�ޤt���4��S���� ����Gˑ���]���,y��pN.� ��9�^W�S�*���d�yuz{��(��hE�Zs&�:�(�^�	�:�}��D �r(�:����Ψ���� ��XD�_��|��������#��xvq�r����~��$�!�ʷ9,Q4ax���:q�Lj��F���[/�����NC�[B��J�m�iS�ȵ���c���.��rI���IY>���ES�j3N7��kCb?e�J�2�p0�<���ah&8�ٳ(G -�%t�0��w�}2߼<e��5��$\ϕ�2�/	�XF��<-�=����^*	G�tB�3@6ҏpb���{^f��Gٳ�z���']κ��Z�d%��p� ��xf��G���gL��"H��S�#@r7�;�RT4wkt�`��/�?jB�	/;���=Bg��>����!�T���W�7��M�L�S9�T:Ff�v<}���sv��Ӿ���_�ģ���'ox"9�8C��%�������+��e�kġVH�J������/�����R拜a��u�#`�VrC���@Z\�lw������1k�����/�G�6wЌy���Ԡ��ThR�?��ݠ����� '�?:�9�pHc_\d�L��b�@�'�hEqn�x�=_�՚@��b��~nZ��:�� �.dq o��?�|�y'
�G�a���ݗ
���;C=� ���;���B�(Q`��E-��E���5��$�A���v�8#��0�̪~��9�-M2��m�{�#& �b���3 ��������D���d� �6�*i�c%�G!���c�-��£|��52zK�QLQ���1�)�65�U�5,#]5l�a<�t�qx����A��R����`�5���s)�j0h�;3���N�?�f[��Sr����^i�O/��_v�&����mgVN�z4��a�U��8q=wO��$��?�N�~��!�c=!�A>��/_��ߊA�41[�l����2�a�1�T��<Y䋧]v(�γc�Rn���+p�QM�4o)w�"��~k���&)�N�/��Ư.F�(>��In�Y�^���kk�Nt�t�z��m�M�O�=*[Z� �k�s��9�;���ݳ}��������^r��f��Sv�T�|ѳב��(w=t� 6�ʤ��̏A׸ۈ�Ys?X�~��NC[�qS�j�^g��zn�_�.Z�]���yU��$�aWu�A"Y�y���gD�C �LV�"՘���S޸4}����>w? �! ,��/�Z����C�Y�~2�mPc��&��ܕ#���LF�ߎ�2o�KGf�>a��͞(4v�p�Nɽ� ȑ��?SBpJG����"��1�]�k{�-7jtE�M�Lpx�[��1�7�8�G� Գ�;�����iI������66a�H�{��K y�M�ґX}D��^<)�*���u-��~2��ˮ�v8@§.YcpE�_>�w��>�.mF��I�g{t7i���.�6����|<e�E�UӔ3E/�W��=
,��Dũ�u�B��wP0�,W-�Ǫ�j>p�lWD�d(i�)�����M�������;��Mrz�^(�����g�/�����#��XF(����{�{0��teň0V����ESX^���|ٱ�H�׶k�ɮ��f�7d��bx{�y|.(�c,6��x�����c|З|0r{-�87Y��wH7+��'�:#�>I�����7�[|Q��2�����il���J�/�!��R���5�z�X�)�fNw5�e��ݽOA��.�Q4��d�W�ΘI-s�y�O/l�W����PɖY-(?�CË���4���Τ(J�?�W"��m�B ����.� 46�#���U�&�����8�Ia�#�i�����EJD�5�wH�2�o�$� ˡղl��S�	*1�Ϩ�26:��"�/�њ�ay�E)f��}A!zj°-R�m�玼Ե� ҥhJ>����Ef��z3]݈П
Ѯ*\n�G������	��)i�h�D1 ���4��2�#{DHU����^�}�R"��*A�@n���!eņE��Z�):�ո��P�=�D�3+:E��Nn��Ļj4�E�G��d�u�0i_;N�����3��}��;a7�,�qU�d��㙨�|�;�JL�?W�������W�Mᵬ����E���/��e�nT���f!�oEj�=!�6��g��s,4����[���w���bІLǰx7ގ &f�8��a��)��M0ф6k=�;ڣL}%���.��	��7�#�g(�]_�-��NF��P�
��)|��n�U׀���=�=��n`��&������
$<�Bô��	bK`��L,s���\3�VK�qޠ�k������1^\E�;���t�4�,݁JZח���s_D��.g�x�/���l��|)�5��Q>���8��e��E�UK�l��R
g�}�o�`��N7�ט�9���_�u\WXO���M�dP��Y�.̍I���h�"��_�<F�M0
v��:��gД����?�=ﶁ��1��:�n��Vѐ�D���BG�$j����"�Q��LN�r��b�:s�/=*~r��peiӛ�G~�1�`�pop3*���jp���o-���Y�5G��6�Z|M��J��Cm1��)�`���o��J-���g��m�pl�yjQ-3��c����zTj�3�kh!�e���1���r��6�|�
��$�^�lA�)��;���˵�&A[�t��I�K}n�������]��@m��i��<�U�>@ۓh�IE�I�9�_��V|>�뽬l����B���Bm����]���h�=������މw��ג�G�=��b'0�\�bQ�{�Wa�g�1�-Κdx-��P'u�h�
���v��3E-#����t�m$��B��r���S�Q�Aof�����p�
(i�$u�-xK�G�6�^��i��9�c)���Ƈ�����b�nz�F�)w�CWj�k�G*F6t���H
�x��V�6��Bc�bq����k���\�DV�K��8�`K�4�!�����|	�jQ�#�"�cK2twnj��l�cq�p�4/)�MY�6�=BO���R��Ql�Ou��e	�z҄�B�8T�i���6��EL��|+4������jw+���Q�,lb��T ��ڽ���3�t2��SO���g2�se��䦵*�I�J�9�����L��d��L�cz��\���:P�5�}J�����}.pk�vBH����ǝ�T���Ҏ�D��y��j�}Sd/Nx~͔҈�9k���_]Ŕ}E�|��O�C��^�!2�6����� %�KYi�|O��ۻ��+o%�dҿn��v���&oCI���~�  ���8��F��"K<A/�c�����5�ge�⊶NPv{���T՘�}E:`�}��閈���B��`���5C�ZK� �G{n���w��`�� G�W�ِ*¶��񠎾p8�aU��������������Xm��&<L[�bEI���bd &º�3��N#���/�{�^J��{�Ms��>��#���$��Ԥ �������Z�٣����hZgϕ���u�k� �P3���I�^0����aMMl�V;ԥ�h���g~�K�5����2<E�����qwQP�yK}�I����8}�a�u'^�ֲ*@�Ԍ��5�r(�'�Fۏ�����Bh���ګr�s2?hM[��}����]j�&y��� 'S0T"��?U;�\D���5Bߝ��ObL�p�ov����K���8q�UrWi�:�92Y��3�@|�(/�6����v�\�N�,J(�����[���z��
�a04xԞ;Z��}c|�Ј��آ�xA8J�IF�ǒ�?�C��-*���_`���'�h��̿ee�{sY�Y}��5s�n�k�,)Qd�|����m��}g��>�cjx�����#gUɡ�}������f��.�M�꒏���x��*~mI�x�tĥ�;���Q���L�滍��!觩,Cl-'��I�/�x9u��	���-�{�Y����sR���L�P@l��e$��8���%p=�Lӎ
 !X�qPX1��9��︜�����ӱ]%.̫�.i�L��mT*�ꋷ��Mx����4;Q�����{"J�L�/ҏ�Z�bּ�K<&�\��q~�3sJ3���.z�m�[*���`Pԭ�ǣ��ɽD�M�>EG� >��y9t�9�h��lȎ.�R�����	��:��%s�$
"��3�7������a�����|Ol	�',���x�5��[=��+���":p{��<�Fp�B4���F�ǔC	�j
��yL(.L���uR�r� �g�HBEM��M�Z�6,L`���od��w�Fz�.S�H����q�2N�J	�R�5�C *#ny��1�W�ǧ,zL��מ�$����8{ls�|�^���op�O�w����g�ؖ��D5�9楞"�js?�˘0QcV��_N��[�b��b�*Qݥg���'�<J��&}�� ���/ ����+�'��@�ϼ�G��IU�KR��CX�L�tR�B�.k�ҧ[1ja���!���ڊ�f�|���7�ȕ���@؆rM�Z"�B:��f#E[�5��Ç����<��8��h������xk>�a��J���V��7��(F��&�0'5�u0;�y1ca�ޚJ��l��8u��G�=
��0�ԕ29�M�=�H+�܇�=3�u��.���*f!��[ǽR�Gi���,X��0��Ùd���6��ާ�8"� �U�,>����-�ov���C���C�����aCթ�P�;�b� �g����1�Ԡ}Ti�+0�G���.̫'-_�9�^��s��|�*|�1�|�4����!�:'��OK�'��ᱭ��!��-���ك��e��6��l=��}%���+B��Qϝh�=|>m��{j,7��7�t`��!h03��
\?�[�DV�o��ɻ�"����yb�ȾYj@Nrt3LEA�	��s�'PX� �����I�e�������3 �D�*%Y���	�DhZ^�Ć2�l��� ��5�Z�Q���F�Y��G=7c���Sx��+2P%=��(��/IZ���(��8������?�p���P��m`/x!��x8��$ �ovuB-�X�{�����M�7�T�Z���К�/к�Ĺǝ��p�f�[C���p�s�R-�j������3��_���a=sO���i(E��"-= 2!u�B�<�D?$�Z���R<�s�v ?���Fo�b�*>��ù$d��  �}����:f ��]�m����< ���rMe�?�JG�R�l��a��}Ƞ��0Uk��CѡԵ ��)5ɝ��a�m��Q�s�]���3G����+�In9;�X��Yu�=���I�:�+��
"?�h�E�g��A����3���Ԯ�|���S����2r�i��x�$��y�jQ�ty i��R`͜�V1T|�z&����]��AɚK�����@�^���Z�������)�\!��A�9���v�{�9yOE3ny��E�
r�����M��즧�6�ߞ_�Q�yRvc�Z}�uYfҧozf���a��<KT�^\���h���ĕ��VB�+��U�f4ɓ��	�H;O��7?�A�Z��+>��>IL$3�;\T]������8I�����u�l��|/[4)7�G�2}|�*�����i�sd@���=�'8�K��];kr�!���U"4nIK_ӛw�Y���:}�^��e5E�.�Ig�,�5� �s�R�c%� �шU��)h(J���V�>Q�$Q|J8�DRd�� ;1�j�_1gĻ���p��`���F�y��mfOYatL��P���b��s�U�0-���C����s��K�[R��J��)l�5�ÊK)��{�k���IE �CŖ�B �7��է���]��m>N�9��R�se��2�K~{�ڢPD�(�CU��<?*Y�tc���\}���a�<R�Nf�Ϭ��\B����u��J�GA4!�� H�<�sS6Q�~0�����d%�\��p�0G��j%�Ѕ�GJ�p�y�Js�i;Q�_@֊������x���ho�U��j�<C~�U����`1�
ki������n���F�7����<wy:D"!Y�_��l8E�Z,�����}$E8��Z܅�n�O��'8��x;z�/|��e��r�0�lo,b)�[�xe^���F,��Ǚ�aH�gq<��CP����R'f*���lx�.�
��߱sp@����_B�h��Tw�h]�4�b(щ,Xw�gp�ke�Dܛ�@�ŗ�BEͯ��Hy�Q�D(R��]���k
���=Z�D�� ��k��eէ�,"��j��1.��5u�o��f$���L����O�m S�'�K[��C��p.x�����2�r���0�F}�3f����q�οT2^�n:0;B+���h����K����L�=�$w ,u�F��2��r�/�������e�L���O�oJ+K���G�a����1� �U8��c70��ż(�˸�f�vp�5\0>=�|�˝�Bօ�V�f�QZ�~�Dw�?(��ԁ4���:zGV�^D�>�JU��F�%ӻ?�yn�C�ƨ)��NEǅ �F�乣���*)@��
�a(�˿���~��ײ��܇���TN�7t�Ɋ�9�'��!�46}���e{워�-4�#�⻥�u����m���q����~#�@w�7R`x�4U:UE;'�T�ր�L�l���bO.T%"nl�LpH
p �5CXz���ʎ����U�oٻydszۦ��mX6=t7�摀SA \ENe�$�8O�`[+LYV��"��De��eSh��9/ 6���{��ɞU������+���MTK4�9�2�{������ZK���ι���<%%����Y��^�@"����)O�f�+_	(�b�l�㡢M��@�@�ڸ��x ���Ǔh�mjZ}�	2R��O�)�m^T<綪��=����A���@��q�D�o0I�A���9k��4���T �x�������4<���i7�qe�����T�9�������lƩ�Xr�F���Z� !^cu��s��%^̠QK�����%Oq`a��+(���Z���4��b�շh���q�C���/���mJ��Anh�uK�^�g�u%5u�j���<W�	*S'*��O0�Q�K_EװĿȲn�fYo������ ?G�q���W� �KB��$Yե_+�D.�$*3M�:��pL�2�H�u�K���B-����B����ڠ�5��Ej�.*����8CJe�˭����'��[�{��D��2�:rfB����b2%;$f�T3W�I�<ͯ�'K?ZQ�[��(����22�w��Q��~݉�[+RO�C�䒦�"=�L΅�#5��G6��V%�=�,���|���K��=���i�h/������,����@�^���(���'j)�35%b]�)ą��/�ͨ���\���Kv�)�������d��
["��m��&m���"qoV�`.�=��t���#�&�)�W%�9�G�L�؋0�<+��Y��xiܵ����x^�!�~���I� �UC��f�AdwTD&�
"���)�ӏ�����n����JS�	3�_롋ǰ�"߮}�c����D�t���8�U�ܡ��a*�c��KM���X�%]s�@��'�"+A��{f��vv^<���]���h��j:Y�4Az�E�#"8�C���Juh;�y`-a��jO0_a,ݰׇ�c�p��Ӥ����AӉշqv8��+�L�jɎ��1�CKU6W5�z��-lӇ�b����V���+��0�W���3r�EпX��e���M'}���{��?���/�t)Ѻ�|�Hg]~nzfxS�tM���r�WC5�2C��_��/���$���</)��4Ѝb��z�7�5�q!���01]�v���I�JQ�\V�
�CM2��1�2�`��(`��*�oY�K��x�/�������U@#��!ݟE�z]]�Y{�������-�p1��f�Nn�T=t�-��<6Hb��^2�n�n&�Y�8���~mk:j�+�����LG`lMR�1�,l����	��I���S��Q�����97x��?�g���tA�i�ۓ� hR�\ԡ�ե0Ӌ�,:-[Q���)l�c<A�*T��ϫ�u�0I#�^jI����@z��Ape��dh��M T�eޫ�����̚���i��c�+Q/�Fm�%z�I{C�C�,$���j�����W��]ܸ5��nx����[���!��>�k:Dg�a�m�B9�zWF|�@ۯUߪ����/]��'1m7%��l�R�$	���@O�鋏�x��ף����R7P�)��-8���~����u��(�"�'�Z��`��cM�[�ߎ���>.}k�Ϊi/�Uۤ$���4ۛo�L/�Pq��[��"�=�̯��BS(H`I��#X�����k�)/�\���U4���U��\��_�D�����2qr�
�E�:P�i&F�/!�������-�@��ē��Jmث@�J��FbJ��	\4j�R�8�����TT�YϢ�;c~��Ӑ�;���Y�s��s�����]"�����tD1�}��Q\�4"���[U0�S9`S��b`��ׄ�]�vQ�k+j�t4s���%yō>� n����#��gx$nr��;�5S3*��)��%gr	"ׁ�`��X����:�[�?�����N��[��f�rS��D{_}�F�Я��(� �SD�|��3���� �:�����x-����e9�2��k�d��/��.� �4]�ӛ�RG��wc\ɇݏ%p���J谘�d�Pq�ʓ������1�â_�؄!e�>��vO�ŝ��Zי�L+������Itz�
������R��? ����R�\��0ɭ�5�~e7�p��m�ҫ��$��S,�x�wb������n+i�+Y��C�w@����&��jc�xBGm��R7C�����g���A���y�U%��1#�ʌS�䚗�y���N�K���@�����^���˛vX�=̞�l!Fz�9Ӧ �D����H�����:4Eq��QR�3��D�	�FU}q6�=3Y�0�4���|v��E��.����[5���h�	�7KE9���0��� E=9C��~ۀ�IJ�E'\x�n���ʁ�Y-ڴ����X F@�5�'9�)d=��fG%�
2䩡M ~갠���f���߃	 ��1�~�dѺq
�d�9%Ff�7y򽪙���xE�j��q%���A��ǡh�f�lg��²Q�%�ꭈ�j~K��A��?�E2�M����`C�RhA xq6��Ax�N���M~i���!p��&�f<�.�x#:54h|��b���N9a�6(�愨|O�鳎2緉�d��Y0I�/�/�W1���ͨ�#]�"S�@ħ�R>�����m�^O�\�˿��ג��c����=k�G��v�I�YJ�}u�?��'5��	~�lj���n |�.W4�n���P�z�ƑFEZ[b���GiqخK<q`�� �x�H��-=Y��ۣؠgQ�VA���uJ�x;�<�M��ao��V�ҨX 1��  t.��S1�Gz,��Ov�T�M5��x�栘��X_>E(yp������,E<`��#�J(h3^�d:�M��ڲ,�h�`�E�~��=N��"V�m��5g��2��X�����G;�F�?�8��e���e�E��>i��Z�*��y���I;�!E��5��V�Z����/=�Zړ�Ĵ���ƏI�Z��h��se�)�ʣLYݳcX�����k��t����?�nЪ���lU?а�56aֹ7���%j�\D�Jl57!ϝ5��GK{��\�t�\�������@�T��_���y9B
���ac��HW�-�W���r�u�̬	~���[����T*jI�$K�1�0���� ����]�w"�����t>�T�	tx4Gǃ1ܔ'�L�|E\��<�N��>s�[P�=��t�������r�S3,��I�D��A��s��ݭ?"u�Hy�m�ѡ�F�ل6ٺ��uG+ e�Q�Ĕ�bS�/�e:ˏ%I�L�*E�_�����24�¿� ^"��3��V��N�w�Yׄ�y���B+Y}V8�yy����tB�Z{nP��苾�aP����~���(w�a_&�Yy��T�/��1��˾Mc'~wb4wܛ��|WY�>�l�N{*R������M�ژ��ʏ���م-�����]�#8�<����Y%�n��sS�XT����q*�`��8�r.t+�}��(�=�$7ο��K�k&z_���P��lhV��}l ]Fj5���s�CJ�f�E�v�:ӧ��哕�F�Y��\�%���([ =�}�R�AJK7TK��G�fiT�i>��DSԊ��(�{����Fv$a[1����c�P�E����D����`6�v��(�c��q�{T����UhO��Aq����Fm�>�ئh9H��5���靄y'���V,��/?.�{���{+���L�?{Qd����&�#k��˖m/o��T�{�*7睭bkHz|�*�݆���w��6w����c�`�!K�D����-�F���e}_�e&�!�
����xdd�P���b�>�_'�.�G1xz���e�h Ͷ��Tp4!$�
2��
Jkd�j��_���U������۝����6�!JS��q}v�����C�[�z�3�K���JÛP!��1���?x������G؋���QT�Xȑk��kv ����$]���S]���;p�?�Z�ɻ<��#Y��|V緰���k�)<����p[�(I'�,��H�[}qζ/�$7֖M�Y��q5h)BF'���} �uXIwЬ�-I��DF�\�=G=h(l�����:��iy��SL�R�s�!ن���O�'���K~���Yb�h�zO�r�o�͍=K+�j�?e��89I�[�׋��%6%lN	�A��Q��8��Gf,f~��֡�̥�f�.��45�K-I��T�>��m�w�Ɩ'Z���� ~�[�>B`����Z���!�����g�v杇�����b;��nj=����ٰ�Y+�љ9�����O&xb�69ڑE���r��k]Ͻ~��A�4z?ã|?�^�(�߶YNE��{�	 �xCE�_�/a���T>�xQ(�L 멫�[���'*B�o�V�)���S�Hdg_5���yÈ
�������z�7(����R	��z�t��.���r�Q�<�����V�9wE�Ѳ_��t��V�s�D��㱀VpoB�6�(�~'R��T�Ft�b ���F�3�{g&������ۍ�̓Q@C7��y�d�=Wt�x�����[�2�hy`{��Yϒ�SY�L�J/�,�k��}֭�	v���� �I�z�'��ZG��9V8� ��Y��[�ʢy��y�r����w3����ȷ�⥰�<�E��Յ^R%x�E���
�KЂ��Em�g��?�X��*�g��Es�ѹ�	%��U�������N�V�BO�N��y�ymX�9V{	��jW���L�E���;#���䄟�Ìr�W��B�Z&�~zG�o�s��n���,���V��H]�C��y�&�JI�R�S����9��&����ra4�/��Ӄe��z��v���:�����h�,	d��UX����kڒttg��~���:hK9h�B��b�jeņ`_���wƴ�7�:5x�^V�ﮔ���	��B}P��@��7�5�8|1�5�*�tm�:��[r������](���e��g�d7^�k8#��E�W4���X�tX#�����[V�ּ�Tn�=�
�m`>�Z���dO�+�}��(/�J7	x�f(�]-�p�8�~�$��+mł<3a��� oaT+��4����sR��� 6�b��r�'b�F[Nt_�'����mm^�{��>=p�t't�1���<�5�p��`�7[ ��C�w�I��t`���|��kk��-�6BJ�3*��tt������~�lw;�rVXy�JR�V|���Ф���eڋaP��,P�bN�-��xJR�ǣ+�|Ui����SU�f�z��@��e)�3�q��l@b�� �? ]�آ|�k[Zӯ��Pn����G8�j��ǩ_�<ܬ�g��FT�8Yh���M09/�<6���X��XTgr��^�Q:� �1��fk :�d��빉��G�Pc;�[�~���0,�#j?���hig���b�]d���y��=�;��V�N��&�AH?G��68OD�`Z:��]��Ӳ�}�:�J>4W3<���m�|>����Y���?���_&V���ܷ�'�����{�V�	��Gl#�a����>qݕi���t�r�P L#�v�#��������1�H��*^�w���ƞ�nz��9��
 5	���S�0�MR+�b�kg�kP����b�]U��	�'�^�6vi'��!� 2]��0��n�}��d�h�'³��@��9}y��C@w���=���@�AC��������{��\����I�����9TI��22ei�a���'�$Wcp]z�Sf�zYa��5�?��Uz���{vL���j3�����M9�W�z��D��i�ֈ��\��N��|��S��s�S(}Be�'��r���ܑ5��� R�{"��z�1���Y�}�,��{t�'��DO	�ުK����Ԙ[S�W�k��bDGr���&ƽ���Z<��e�oT'��`����C{������^�rcFoF���Ϫ �S1�(f�Mצ���u�OIg��%�{�A)�����_�G��>OX:�=$U���Q̷��S�*x�4�y�(������)-�;V�b�<��
 a8.֤��'z2-?����-WY�J�3nTfɒS�i3��.4��1yߍ�\�5mɝ�`ZC[��v�4��o��/�%��I6�v���l��?����]AS��踇]��2�Ц�{�d��"�`��v���#X�fK�Yw#��x�,�
b!�|14(M{���ZL�U=�]��WV�t�p('���/����k
������6��/η�^9;�Vjhw�"_Dd�xª�_<Ҥ��r�0��B�ꫫj?�9q�!���@�
�c�f�;+��v����� �{|\o���br��6��)�D}Y�S��K҅%�7)?c�?�j}ط*Ag";F�ơ	06����@��;Iy���Vt;h�t3��xƹ�#�C[o�������s��6��H����P�B�HW_�����3@���
�CR��.�8"W*�E�(3;�<�`v��f�(�| %�,yQ�b��z���Dl�(��a��:g�}�3��-׳/VX4�M8ծ���Ȁݞ���%d][�N!Ε��e_wݢ�t����-_	�:��Ε��P�3�'���6�%_r�M�5S���n&M���ϼ�?e��x�k�p���N_\��,��;�A���iK)v�q�5U �&�h?m"L�S��Ku�}B%a���
��9Su����n⼨�OL_�}���(���j��6ÔXO�!G*2I.Rq����� aȦw�(e����<�7E�!����aT;�]�pfV8Ͼ��(WҔ��#M����;Ѯ�2��&�}��:�k3T���3G�7؈|�w���,��o�J����Lx{dmz@n�K�����þ�̰:<����e���r�W��H6#�����N�����٤'r|���`ƷX��'�z�}R� ꠖ��Q*�q���]��T����-'6���f��2�]��w�� ���pK(G�V���"�����9{@�[��Z
'M�фT��s��l�?G�wf��<ꨁ|0�l���(��i  �BΕs��uaG���/���
l�x�`�oi��	R�NY���T��Z��$��W���;�Fh��z���� �bY��[�L�
;u��uܳmh�3�t�U1;ԯ���aC�qs�EFó���0�i�4�׳�GM�k�_��� �M��{�m��
���ZN�H�J�����L�UZ��K�� i���COg��7JL��k�������Dw8�[RZ���,�/yg�T���GnՒ��-#C�@��K�����ǜicrq^�J�H�H�,��c@跀,��A7�4R���gLXؗ����E�uil��'��ne�e��zyn���ij��];A��p~���;>�b���Nj�+CL�8�Ƚ[���p�Y.ij�ji�*����RTU�r����#Û�Nw�Y��O9~�؇��}�y*�������3i�R���|�}��m[t�#�$�u��	NN�㶸I�R97���r!�)� �|��XA�!��M-&|��w[��]b&��Cq�l \{kC!K�l��N�uQ��{\wj����� q��2֛"KrM',+�Ή2<�?��᥄9l�zd�Wf�<ǸZ2�?�J���>}�j�M�����S��{(��˂�8�G� ����M*���z1Xf�$d.4�e�6�A�7TRä���0��H��G��#r����*�F���x�.���c�O)����a f�ho:b��?�s���K2K�C\М�-!��j����d��z<���(�q����8f-�dEI>�ph ����I
��_�u^ �@��"�۱�y [U�/������e~���ծj�엇�U7A�M��k�6
��FHg�'f�
���(��0��5��l=����'��}.�������/=���;��r��o�$������"EA���ۣ�sw�d cW�x��p%�����K9���J��zq_�2+�V���ˁh�+3lĪfz)�<�C\�	����i�j�[W�ߨ�z�D�E@|e�Z^ߌ_��}�G�}��NE���kQt��2��0߿m��u�2��4��'f��v��L�l��+�Q�]K3>j�p���	Uɫ��E��J¤M�/ù+��w-�q�3��9���V���pD�͌N���;������V��b��y�!��������B�?���8�m
�х0P�ן������*��Cefe
����WQ�� l*�����p6�#82�g�
*�"7b��</�S�ä(K�Y����P���4���t?����۝���v_/8��[��a����zꉺ�au�vw��=���Z��>��f���.r��/(�|(��Dv6#AL�Q<�)��:^=pK̀|�|Oy���
ԎDW'�o���>���OYS`�݆{�����u�h��P8BN `8�Y-_��y��k�s]�m��Q��iv����*1�]q���D��M��7��o�vz$"v��OQ�̦�YEdOITа���j
��:�^C5Z�_�״|�߬"��scz��ѣPJ����Z��̋~�=Ah�_�E�)�b��I�S؋�[G�!XEWS?hy'�t2�y~�x��Χ�6��ڒr�NUv����t�S�����*#UVbT����xj������e{޼�:�d�ucW�Q��-�gc�o+X�� -0�}d��>����ёƻ\p%	�3�����	�'��^)�i���8�T-p�bM���W�L�Ѽ@9�?��[���Y���of�lL�cI�m���@��`�$���"X��>-&��D[����7	�%��Ǒ�o�}F�sY�i7�9-DV5��(7�S�0H��y-��#�
Y�3�)aPA��O_��!"~]-@��!��!:q�r2W���귳����@�A\\. �e���Ǜ��^�k�W�rׂ�@�E)��]%���U�9�O�n�)q�	y����2>;C�;i��;>Ae�������]�p̘��s�{�Lz��kf鈼S ;�&�4��)�D���Ws$Z+˩䁉D����	�>ꪭ�@o��6	����%T�����BW��_Y6�kaWlL�)C_� ûze�B1��XXbx��1}]\S�JR�����֍�Jk(�X'�`���ay���4��0�}>���'��6�tt�;�lE�]�>�	�o��R��G�2�қ�=nk���6c��,���锑�n�j)�>6���E�Ȼ����������$��F�+�v6^���6�BWQ0*�L�@��ȇ��l�0/j���$EgA���y(��c`�M%˙`v��ʳ(�Fb��w����/*|��Gՠ}>P����i��@4�IW�72΅��--X�-���������
��#ͥ�+[��N�d�/@q��MO~�����Y�u7�X�ge
 �)��4�=��1L� g�:��$�-�1�s+��n�xq�(g�y�xd2�J�F�j���S�dQ��q��9��ڡ��3��l8�����/�B��������Fk�K���(2}�~�W�ڡ���I��H4Y\�Ya��a��H��w���ļy���?��/yZE������ �n��gQ�K�9�e;�vﾞ��V�feI��Xϸ-T8i7����d��
�ˀ�t�ĶóKr^��4{��gf�w�fj�t-��ɗh�9�8�J|�o�|$P��ݘ
C����������
i�����؄]p��b|Te�+YX��4�E��zv����H���K?0>���s�ˌ��s.����/@�cQa]+ȍy�` ��69�G��vc����Kh�9����=+Cv�.��ȃ6R�O��F�C���Ɛ^��;��<?��Ň�t7�����8��O�+�$V�����n�B���K��z/�Y�����ȿЕ����r��l����5�am�50��K���oh4-]`�O��K=^;�ڼ�kܵ�b��۔P��R$����G���vg%~�~��bja~�x�+�&X+�X���M�^�Lv�wy�X>-泖��B�nJfiQ�&�;�|1�d���n��62��I�C����)�m��:�o�~�564����w$�$&�6�u~��,rk�c��R���}�<��B����<o,S�4�T%�o:�1�3���c]��@�Ո��k�^_�����buu��)��!R���u�r�?��M��*��Au�Ҽ��;�nO���7R���H�*-Z: "��M'��WÎ�� v7,k�� ���ɡAT��?�@��x�|*��6��Z�
;��b�c���PS`ec(s��9|���=V�J�7+ܛ��s�i<�h����K��+�㎬�)[��tD;���l��ʚ�3�sN	%Ѝ[�p�Ia����z|ė�˴i�Kx�^���$��l�>0H���}b��Lj�l��F����+��Q.s�4�!$�����P��o��E!��C�SH��j�����jX�SQ��^�-_����Qh5<��i�V�x�J� ����P�'^$���h��!�������Sݵ��L�ۚo�ؓ	���Hx��\�ǵ͌^�%]W�<����r���9?@��2��ٵ̕pwy5`���"��M�/��.}��uA2!�[#$<͐b�~:o�y	����XYvP��!D��v���Y��$,�,l����9�$l	����ܻ�)b��G�p���M\`�'_f��m2�Qe�(U�(:�2&��Z0㢿)�����}����{�����2��(�n
>�)��L�6G��#�i�~���8�Er�)➴x3���?��C~/58[�������h�1&rO�g�5ª��%��	j�'Ao�^��±\Fw�oP�]k� s\x��0�vi���W��y�%?�8E�l%S]Px������x�L�˽D����ч��T~��NM˒�X#E��)���)����6�'k �j��=�X��RgAy�Ä��fϪO��I�0�%�W-��c�� ��,�1�ȰˬwE�XGs~97��7�Q���6�;޾g�g{��&�1���H�(X��sF��C��G�|��bGEr����!#��:�S�S4xDy>KG��l�����X7��b��[p�x۷@[�|.na�����Yh/W8LX���ߚ)�,�t�>@� Z�}� �����TP��əd��>:8��:���b�`����&׍�}�w/���]][�'탢�Ĵ�q,�Ϡ�>�]`e��ݻ_r���יڠ�b�����Ԭ�C"�)��!���G:T���) �  ւbI� �9���2�'D
BH��B�f+ hI�[��'�[ff��YD��1MYǩ������71���p��*��7��6�{t��:9:{|+~�p�4�1Gc�0�n�J����b|>b}�Ev�\�"�xKI�8���T[02N����0J�X01�۝iU�|�ֳ����-4��P���%����⌿��9٧�'kU�ue�];�Mb$�m$|!�]=���Y�,]0�\�䖂��5�����iNLE���H��E- C�������P���q���
f�m} ӆ��w`*վ���&k$>���V{ٕq�EQ�1i����v�� 2�)�ռ���!�pmA+�9T,���M�AK/S�_@��v�:����ﮔ(Y�%�ۤbY�K: �U�!�l�Yx�}H?�,��
g;\~9����D��xL濾�	�3���vz��c����Rx��h�#d4�8��1`��_3��i�|��V3T�����d���e�K�퉕�=wz��%R��R/�E`���f������yFu\�}��v�ɒ��S� �Yv*E��qߥ}�Pud�a��H��Pw?M24ɏ�?�Ћ#�S����C}fq�ML����z0���Ef���R6����8�0Ĵ����:d[�F���u��Vpx�B;Z�HŬ�R1c1J��Fz	e��-�s��}dn����#�5��|��h�<�X�������4ۍ2���lF����
Hi��)]M�f��)���ǽ3l�˲g "�t���H�\.F���_�'�S承�#dB�Z���z�����8��`O�e���Ւ!���d��N"� ���L��A�]s�x��� �����pz�9!]w�Y��h�C.$#�\�gJ�x������ �p ҅hR�k?n�I�;'v�؟�d#m��
@W12_�D�[��U���"��o2F��1C��?���$i�k`� |MM
�y���>A�Oufn��`�j�b����%љ�M���͞8�����ۢ�}h�i�;��2/�٩( ��@��`FanslFxF�Qt�|u�������(�熦}
��PI�5/��6�#[��BG��{�[���c�5�ua0s��k�����)���9���~�)V�|�q�=�6�3��pfD��$|X� �p�g{o�㑃�B��/�ڇ�6=��_�W^�NK}�.Fe'?tH��M�8��#wd�����y��Z��Y(	���n	���(ߖ�a�N�bW�d�S{$�+����ƀ3�F�N�P7���4�q��_{~��)�/Nr���x�Im/�&��r3������W���H(C����GP���>~��N!��k�\��р�RxA��K�~��abٶc y�V��P(��[��d��ҨG*@"p�W��tc�I��+�`Q'��zv2�Hf�ci%i�����ƛ���n��r*�ꬢ?1�[Ǫ0��`I>#��(�r����_?${l�a���&�y �֐���q5�i�I}���D��T�O2<t�ķ7uo0�e2�9��"C�nxim��|T\�d"@He)"oD����{�~2/ɜ��6B�ؕ�,0�8i:��w�6�����_љ^ǼpNq�
MD��M�B�f5�b��������D�)��Yv偅N��"�Y�Q�K�Vr,�@�7x/���b|���Ȭ-6D*ҽ���*�%���^�h�r�^�z���K�:UI�w�-�$�;����M'����mi�����7�~.]���;U7 ���4X�����T���ԏ�����&jY#���^��\��r�ܹ�����[�kh
k�x���/��
�j%W��P��2�zb������#�Lorp���[uϵ�;���O��Z96���Ž1?�	P�Ť��T�x���a_�p�MXgR(Wd��`�T���I�z:�=R�� ����qٖ/c�����*}�d������{@>y���p�< "_��=�c��㽥�����+����-o��x�S���9�M/��a��&�0~WG����1h�Q�Ɂ"O�I���n��HE@�>�.)��-5������WN�~;�ǯ�<�n�P��w��K�pbr�7�� ��=0�'�5��[���-ںCl��[�j��N�]�#�����������׽g�׏�҂)��=����;���j�Y�Q�۳L�	��0oūɄ����P~�HM����#!_(c2��,�{Æt��1��Q�_p���^W�K�.׀ʜ��F?�>�p��&�g�x��>r wᯉb�EaɱԵ;�k��+`�a��Z�ԧNr��$p�pk�5��-����ĎҋD�r�&;�Z�ҩ�:1��X�ɒV�OU笔�w�f�ܭ}7{v����;Y�!y/[o�_E܍Q%�<H�&����g�Ф���#�J]�N�j*.mn�w��T��I��Y��yq��^�L�so����e���|��;���{�Ҟ���������($ujW�Hh���Uu��a�ĵX���=��$��K�j�L�D��z�&�7�wH�-?*0�wY?e��
4�s@t�5�m6q�bE��O.�e,F���.c� UK������-���69����́D����޹�AY��*�<���K�#�z���Tz@��	%�pU֡Z�I��^.4�3↼�?���ԧ4p�3��ǿFTy���0gb�fӻ���-[s�g���#m�\TS/rYBrcz�U����G"{[&��sx�%jÛ�u5���p���3��MI�
R.��B��QK*�N~΅�d�8�U���[�v���r�mIq}qA}��fD�4J"�,ҝX\Y�Z3�$�wr��iI���&
�X��vt�.�F�a;"��;ck����O{C����965]"Q�H��p@��;�`�y��*����w߇�\�$�{B����p�8�uZ&��]�t�+V̀{Ԗ�w���UMB�9�27�z���E'D���u,J��o&��q��!��>���e� ޿e���!�C:��j�9ID�S�í����~�x.a�
�X�b�XR��S!d���w�,���{��{]\�n>mۄ�0m�3}S]Ց^�I�[�!�*q���_Bt2�6�x��
7森�L���*/^o
ve�����Q�io)�G�a��XV�
�C�l��Y�;�g��!G03?����Қ���EzGJ/�i`�[8�ʠQ��|:�A
���Ȣ��k�6��'��4]���2�t3�L��G��6��ba�x����}2���y�~6��K"��l�=Z�L-)�[>R�8�S��s�<̓6�̤<�¸�ע'q�[�9�'�!�uUN�A��4'��@VC���(T����f��|�C̑��RB{G�`�S[o�����/��0�m�ħsMh�g}Ih'���>���?����E�Wc��g���o�m$|
�7C���ϴ���i/�� A��Q�>V2F�-b�wGR���������N�VM��ΟYY��+Bt��'������n-��{�#���٦_Ў���Mc˸[��������XR:�51쩊W�)���\ʏ������5e`	�^��/ I�u�]����9 !�������V�H�9�����&�U�L`>����7�8�'2t�"J��2�!$���7��3�m��>�-f�'��O�m�V�(L����RKQ�Rk�Zn�~��*�?�-�vK�� f�L���T�◅�1��}���7c��H�����$u�m'��.�ة8�{U�@��Q-����>��z�zW�©��I{�}�g?�Z&^8�;�% {E(����)��}JX�Cd��~L�Z��,�|��B�/���r�I!r�x�}��S��wK��YT���"��.��ZFL��N�2w�I&!��B�7��^9�k����8R�=ɇ��|�'	�S�w#�6��FP�t�R֥ӟF ��#�υ���!%�H~�l�ac�������F��B��G%��H֓fZV�Y���Z�TuX}E����i�M�e�B�q�=�(��c�J
+_��z�S��O�	aG�w>Dp�h�嶗��ڜl�9�Ml�j��S��$��T7a��٧��Ǭ����,��w1���*���񙥅�`�9:a�E��DZ��a�0Y ��1��K�S�\��̰M�e�Pw/�Z��]�A�V� z�^H�"�@������x�:Kqᄡ�&��S<|0V�F�H�8��y�Y�Z�B���d���B\�z�L�\9
�K'&�xQ끡�������x		.�H���=L�� >�'�����SY�d��D��z���2d3J,4���>J����i��Ib'"�z���>��˺� ��P}����q�y��V�������S�~K�G�i�j.`����蒊�G�"S��"�F�|
�Z�u���B���Iu������]�ܰ����^�D�=N��5���+X�Ųq*�uw)U�,������O�[c��o�D�&��4Q����V�ɿ��iJ��/5�Ff��A�F�<7w[+��2X\·� &{���8ᩑ�t&��&#;�,��C*�P��6��~��( E�&���",����󳃢�}#E��
��4�����8&*��Cp	���
s�`!143/�/X~~-�B{����6��i�b�?|#�����7K���Y�&��M�q��P�M����\i�����_R������h$�Xm���?��Sͪ� rЀ����c���6�<�|��]KY|C�U�+�#�Ǣ�s��@߶į|{��!k	���U̇l�t;7�������|s�H��`�U�Y�1�t�5�����`6Jc���r�]Ka�֡�%<Y�Wr9�0t������,1���h�X�o�{S�9�f�3�������E�)�:��!7��x��Cxnk$;����I	���bk�>���P;����N]K����SLσeYu!h/,����@����Y�۾S���o��/Xt��h}�x|��V��~78/�F��C��	�G�O�/�t�M���l�}�A���(K4��PS��Y�(�Q6dD�b��˞�DJ�8���@ �d
�YEt�,(ۢ�G�.�D-��lY	�@������˭%�!LS��G�w}7����.�d*��c��j�X>����K�U�d\��oS�e���q��t�ς�@���d?�>��|c�39�V��mu��X�f�N����I?�9�f����[�� qNyD��ϕ���쉦�i]���ɼ�>����AT�<]��o~Ri�Ж#7u\cͺ�~}<���D��q��1{�VJ���v�@�ɜ��S3�\L�R�j���Q���+̓���p=��7C�fPP@��*|�y��K�ot�D����/�,���O��q=����䂁x��
%E���2�E�����7���'�E�����rU���Y;x���q�`��t`�$X������2�B ��@����ov��*�ϳ�vhuWXi�(�>����'l
�V9����fl�K�4��*���L~����P �;;ک���=�kx�Nġ\�s��������O�_T�Zb3҆�+F����k:0_F]��¯�懑`�8A�2����1!t;D�zѣ������->u�Ge�r6��yK�R��g����t�ōR���5���R��,���eCהr�"}�#���ر��b\S�`��C�| fK=1u�����|沄Fty�ho}�\�# ia�8�뛱�T&^�&Zv ���ξ>B��h{�Q�1q�h���
�^C��Re�LC�W��]�����}��ho� ��:�!�&���m�c:c�@)�Ԉ��E���	�W���m��$x��j�?����c�̕��{���S!��9k(����$��S��nہ/�x),�$K�9{smnn|i�7��I�X�y������/�;����x�{��Hݗ��j����V���=�-B���5�O����(?"H?h����+� �YԑҬ��m7c��zx%Q'����F�8:dX�|Cy�.QSY�$Ty��龎M[�؆��bQ=�����Z���$(o{q5�lZGA-��H��F�p�#&;ܹ��n�]Kp����F�1t`���1�4>���Io�z�u�?�Eui��8� .���6��56ҽ;/���ݺ�+D�P��)N��$%��ۆ�c1(i��!/��-�2pw佭�� ��GZ�N��3c4Cn8��`�YT�k}�T ���L5*��k��ƍH�ב���۱��!N0�Z�n��GOΗ܋},mP�?��V]�.�ƹ+ �|�
���8b�_�Hx��^$L�;6W��˱Q<o	�T���~/:"��)�L'�pvd�t���!aTG��s�U���-q�֕�ź��)��#&`[���!�36-�|"�!.;��P[���t��L�߇Y�,�I�We)��k$��|zDt1���A����u�m�Ь�4��nM�;O�G"����R��K�������~���1�#^��f��hU�	¤;���ˡH^�����.�r,��ֶ(H��͈�"��/C�A;��%/Û:�p��Y�����vRC�#烙�Y�f�+�}������!d����Rb�+
�y���v�XN������)���S =;�Cr]����f_�B��6���cZʩ�����0,EBQ��I��.PD�7��d��A�%߷��
�f�>~�]�����؆E�m�z��p+"�Q<�~�e#H��r�nMTG���kl"-j�@�e�+�z��3�}�.DT�K
]w -e��,��}�s�T�_>ρ���Am���٦�P:���n�l<JN�����d%'�:�� ��a$��^vV�G�f�[�s��f����bg��b�z��d�s�$���^��ǈ9�Qc���*K��Q�eQ��m^qQ�HZ��],���
>5WSIk]��z�'<�ʟ�Q`���~�������!�( l�l��¼���%oo�,���?H��N�j��a @��ߡȘ�Ƙy�����r<�⢷�58�E7�bH�t ���g�x#A,�s:��w~����v����_�Z�Xg���ְwø����1��f�+�n��[s�4�.h4hQh=��{O�1�ڪ3u~&�˗��@��b�N�0��2T�b��8��v{��If�pߍa:v؎k��@9����2H���0ش�Hğ����i�u�S�("��Dk(G�E7$I�{���]��NFNU#� ���Y)��'�d2�E�߃�~d�M�\���������i�yզ.����QNj�ݒ�*�Yk��/�l�JM����-Tr���dU�b��
M� H�@�߯^�.���s��
�7�b��2P+dKJ	z葄������v�t��U�g��s��,�@�x�׸2�(��:��wRHԥ��O�ѥ ����J]���L���7ꤑ����??</v���������gD-���R,�[][���������5�hZ,=�yp�c>� PG��x_���}�q�`5��P�����^ {z0�f�fؖ����y�@*~eLt`6LT��u?x�Oɱ�pВkI���  IPP��X'I�F��F:��R�	7�{��-3�b���.��/k�Y�Զw��B	�8��`�)Kr�_��K��]4��*���|>����ƒz�x&v�8�Q����'j45@V�ݧ��'Mc�؆LE�����')��g�i>c�P�̢D�)j<���h�:�6��l�A�<N�����ߏv�#�c�w��Vj>��T?�\��#�A�C�ƴV_�ͥ�D너����"f��p�ջ.���Y���^�Iˀ�#���zqH���/D���t�O�L��#~ݗ��":��">��E/8��5 �??~o�|��b+G�_b�#3�r��lz��r�v;���yQ�'�w-I&�W{B�洣y�s�i�Roȩhk=N�NUi_hT�3j���n��i������V�� ��ʞ�4V��b�������'f鱟|����:�뛓w% eS�ݡ��js�����p'�ke)�W]G��x�m�x_���I��l�ھ���"����<�;Y4�Sk��|K��1����N��º��T\o�	���/e�h��ld�-	��V���2�E�cO,4$������n��Ϙ���W �!\|�R�)F�E �@�ҋ@�0�����Vo�� S6���/?X��Ž�Ù��%���(J��M��R�k�w��{�DH�؞@u����4����Ԍ�g'R ��.�t���/�%�_�ڣrp��D���|�������'\�9��NJB�19���R��P
>�����@ŀ�uz#����#����܈����3���ԧ�h�=4;����Fߔ�\��+�:_^b���gBX=������^_�Yh`*����
u5vL�C�������'#P�PHGU���xĊ����Ǭ��l%!���6tcSL��X�$�sX��@��_ g@%0�Հi��cRV���=��#cEN�LcH�Z����<j���6�޶�����o��h��kz�5�y�,4n���܇�W�g��}8��;���b�ht=хR@kՑ�1AsĮ�B����ha���{�/*�٨�1��g9g�9����r�(�UQP
�I�a| �C3��X����Ma�s���Z]lу�<l�ڒ�W2P��b�ƒ�T<�b�M_�o�G¦?)G��b P�Ȼ&�~�(_Dm��کPHNdy�(<���ɭ/uD��j�-7��Ac~���+HF�x��|�Oc���[1Ϫ�x� �ߵ@����S?hT㫢���-���)R���ێ��gh}��R!ۆ�Vxb�F;xtKE��h�J5�RD���E�Vjv\��x��Ŭ���'i��C*͞�]�*��g���+��n��l�cW�M���n��2D������L�eJX"&�D]����g�����ʹت����>S�Uzc	V<
3����F4�^��g_�G¹�u��A��Yj�k�g�V�j�?X�,��C-������	u���Bv�'Y`5��1Z6ո�9��Kb2 �� 6����1�*��ҚDc��7�B�bP �v�?����ȹ�{�&6�9{���:�� �����0Sw���/lu�0��3�T��U�z2;�^��	���v:�� ,Z��k�Z�F�xYz7U�7mMS?ld�K�V��#sk���'�-�j�e��(����\�4����q�[e�4�a���0�\�^`h������2����"�T~q\����^c�պԛN��×�"aQ���#�4�g�	��j��g�Y���x>�ڐ��z������3mF@��q���RH�Xڠ��M$J=*�	��u�̓�3�5���dk�Yw���8����� �	Y�e�d��A�,��pC�h�Y��"�D �k5����7t ��m>HJ$��λ*�0#i��gx4���
ڕ�Bܥ�\�.B̰��#����%2�qW|��Cq�9��$�N�m@��?+�����`�wt�}��'�B���{���K�6JT�#~`�s�����h�kQ�h� �j�W�`���(bb�y��Y{y+��Vu%�~�[&��e|Aw���,�}����u����X2�qlN���2�rWa����е씶�ff�Ay"�E��!�$�����,� ����Wa�v���{�˥:�es[,���K�v�`ޤ�Y��=�&�p���H�^���.���V)�z�6�~���,�#X��2��x¿��`��ZOM���#���O����d}���iY�O7��N:���N�=���<v�8q }���#6QV�6,5����f��}��PQi΁��:��gdY���$C��{�0w�2�\vH����`u9���27о\P����z'�N%�3;����Zn����,B�K������q{F���<��"`c�g�
�9���]ʳ���;������n���o�0g��Ċ��V 9����h�ʱ��y��RG�/��� +��p:�O�C뢑~�iW��
�|��(����|\�pe'a��(s{�r����Z����&ׇ=>�UtIa��r��>1,�6߯Q��7�q�Մ��A݂�[�r �	�3��$Hi��s�Ry_�n�J=�U��3{A�,F��o������[Б��H��ć��4)+Ȓ�Hz�"�x���e˳�^=pm5x&T*��E��K��Y
P����f�7+�>� ���ϼ:��Q��N�~''ӕIr6:������@?�A�D����Y����a�qjp������Q�" ۾�n|���UŽ}�ڼ�֒�ZG�A;z_�.���Ъ����[�%7Z��f�EH�b�N��Y�jF����&iv��-��G�!��XO;rm]���7�X�;��w��륝���V8�����Qf-A�;�AS�us�B��u�Tv����j0s�;��hPV��Y�0�Q$��]��X�rkoa����ɑ�����* ���K�/U���q!��͒�GOr�-g 1Ux���õ�B��	0����c�+�p�A��������"�_���P�%��L��!1n�U���Q ��m���r*PhAE`����#�;������p�ÔrN������,/I����I��gL$�-7s�Q�u&�P�xH�#�AX�������n����U�'67�N���ap�!�~�b�)���P�ib������+���E�>�sU��������7�R�M�"�ҡ�<㡴仞�͖)^�8�D���Ti#�ր��B�<�5vjq���u?�aQԌՇ~�� ��mK'C�W�u�̫l�SF���`f(��5*{-$!���`�%������#�ڹED/�eȫ/u���%����菦�f�BC�O�X�w} i�\ ��DGa���87�9���=�+��K����!ό;�M=��G�3$E�O�Ft�/�Q͜�e�!�Gl�Q=P�xA�Ft���Ѱ �$&���{���LX��
�+��w}�����_���-��͊�Qs�\�����B(sH�É�$Q�q�6<�H�����6P�sx�nv��*����5y?׶�֢���9� ƍ�1�|xV0J��?�^H&a���1-u��s�"P�Vt-�(º^0��#:9u�X�#{h�0U��β���*��	#qmv�T%R���ݗ5/#�B!/������E�J���m
�"���Y�seG�������҆��6	z`��	��n��v[_�V�0�xb����,w��&�qw�V�b`�l,�T��(���޿k�m�D�;�z�=O���� ^K��-,{�C�.�G�2�ͤΤ���=���{%�1�\��Pr��'.����(���qyVRo������Y���]ŵg�%��Ƽ����ZS��v�����[�C���ɱ���9��å	���-*�J�d��N��"�i�N�љ��������j���	�2�8��0�4��{[���Z�)֋HLM����n!�y�ٚ�K�j괗��2A�@A��%���k����G��b�d�����h���	ԓ�i>EB�^�y�����5�p���y�'��'�ڀ�+q�@?����W�E}�Al�'�>s5�ʝ���W�{4�
����
��%P���>�&K�:�����de�]��a�a�
[�h����i�p;o�e;�l����:����v9k_�V��R@U��f�Hh��;c��Fgb4����(G\Gm�+Və\wA�q��KJ�(�1�76R!����C�=!�9ҫ�J��Ѡ��E{
n#���V]FN筠-����T E:�Iil�@m4q�ov>�D���|?@I�R��z�Y�"��B]W�J�P�\�s��(��J��I��!E�Z4�W�s\�r��.�aJS�?c*��m�:����n�q���=p�ER�z{'9��1N�p)�,-�3 ����hm�jN~L�uh�qҾ`�²w�3 yQ%[J�1O-:0�4Bs�������<���P����[H���ψ�-` �L�/3V��1��T"�{�Ǒ���v��)��$��/H��J�B�'h����Q`��
2�9F����Ҿ˰)XO0壶Ll��c�pj�K�Y�U�7��8N]ug�>�"D+��2~*HW5�����e��J�3�j�e;�LiO6X6��t�7�Hc@T�K=�QOf�w/�ҁ�������� �e*������H=$�Ȍ���W��:n��S�h�v�^.A��S��̢m�ܞX�T�S��$����LA~�MH�	2�\�z�!*�� ���.�ת���ˎ�����C�̢g��A�����)�k 7��z8v����4�A���i�����xl�:P�ǡ��76�Q�'�$(��^W�F�pi��q�:{�-����#�>x�D�z��_ɼ��w�J�v�i!�܌o]OC9��B�;[�~a���L�b��xx�ۖ�.�.����k��k����R#l��W�;��X�rF�N��W<:�ǐ����c�c{�\�FZ�� c��qa�K��o��٨L� ͝GO]�8jD��|���O4�(��si�����ЎW#�M}�p|zI>J�1��	a�*84�� SH��l� 
odGD|a�Pg�0��>�Y;{.��]��a8t�9I�l�q6犥�s�Qp���EX����b�̖�<�+M�ū��씬����`��ƅO�I�O�[N�ٺ�&�o�LL�q����S�G���a�8�g����`�V�*a���0vc�xW�x��������u��Yg|�>H�jk#B���~o�J�AJ:��-�0� ��8\aSr,�b�"Mz4���i��Y�Ӊ�T�MŇ��7�U�%������e���qِ��^a�B����r�D�*�<�R�dtB�c�$;l�s���1�)5	�y%�R������T�{}~k����e�r&]R�����d^x���i�d�?"Ftmv���Û���T�c�g����^_a,���m\Fk��F/1���	�ZZVAIA�:\��z�n#T�a5 -�����j���OlX��6]��|E�˸x֋��sR8ͫ��^�;�qM@�fb��R�	]�iu�y�k�W�IY�W��F5˘�+:n~ĺJ����|�O����$v3��N ��;XPN*kU���r�fup�va�d�gp�� 2�K�����ñ������~��I�P��S�4�D�c�9�/!DY�!��ųO�FG�y�HMo_ix�~-7��{����͟A}߿&��͡��T�W����Y��b܋.��R��օ�}��R��p���y�g��4fB__
�/-T��
�e6'���7cA+��B��;?ƛ��� �	�Y8
��c����(@�����Z��EP�teC�xr��{uyહ�A��N� !�����Q������Zj1��Y�㢔��}�.�� ����,�Ɯ��f<�^���`��T�I2���?[M=�E�=�Jx�)5����cc\�	a1�L+ݢ���=�@6$�G0�dY�pw&ZrQ?�����,u�n/{~��M7�H��|�Jf�������s���ؿ�6,���\h�s��b}fb��t��*�d��T#|���x�\!"B�=!�Q�AG�ϙ	��B��.����W@�&.kl��>�ܬ�x����}}�!1�>�l��c�����
�G�v�%͵�l�ַ1� ��#��a�_B��|4�NY.�7��X��S�Ғ̉��9�2k�X��E˷C��6�\.J����kϛ���BzƐ�\��hI�-_�
�#9��K��U#��f�
k(٬'*;�&�ՋT٫>��������vw��cc���]��%�k� ��=MSNCTWї{ ���ᰓA�� �4���8X��&}F(<g �:W{bN�F�T�
�G|���5:��;�o��6�;�Sp[XO<@3�EL�Jz�4x;�t�#�i�d��O�4g@.��'��� ��ji�_Nc�7N��(\�$C]g@��\#�ҝ݁���%��?��T���/��l{]�k�Y��1�:Kxo���~���Nꎺߪn�
��n@;J.��ݭ,�^���`�_�W�7��P��\UKH%���<Ǟ �?
��*�:YV��[0�;)�.�5:ȮC=f31`~[>XVÕ��J��f�z��j?Q��}9�=|���G#N��.�PaI�N�ڧκ��V3�	{��I+C�D���L��Qm�UI�``Ki�Q��d��� �'�-���fcK�(g�@Z�W՞ACc����O�Lp��:�Q�GX{�jƯ�A$�cu��F���	A���VHˎA�tՆ��2p
4���w�}��mo�MA�$)���XW}� 쿜���#��7�zc{�G����j�C��Y[�	p`6l��w�h�0]�b�6-Ϡ̏��N�-�2�9�ȍ}"][�^ҩ��������e�Z�:T��/-%w��|��G'`{�K��!���$��$Ш��K�j1�8�Yd�.՞�DO�yB�x�,H��ݞ\ڍ��W�zp��Pל��<42~V��-l�}m���w� ���Pβ�@=m;[*$٧`�Q�������YѪ�c.��Iv_���gد�?c��Ou�7���ι>���v��<I���Ph�`-�	u �j���!P�I�[>�Ȏb��M�yp#w��'q�=��� ���ө����I_AF�tWVftPd��k?������?�\?�ֳ�E�R46�3����z�**>*kǠ��kn���k
��,���OઈkTz��3"�wO!ȧ�U!q�!�"8���}]K�nɆ�Z��^{�:lT��;k:�d�3\&N2`�8(��05��li�zv�
���(K#���I=��xm�b��y�V	�2��3��d�-'f��o>z�Z�#��/���I^>��+� O���M�����a��N�J�[ x��	�0���~��x�4�6�y�?eRO��QkТ�<��(X��?�1����e����c�w	i�o�>�����m��@������������wt�/������2��ZaӘl7�t�Qդ2��S$�9=#�ធ�K�߅����0&M�s����Q98�i �N�/�F��A-�	6��6��w~�0���8ɴ6��P��T�Uo���/m���:�V�*2y�6`�����v�c���x53K�m*�b��$~��*�ȢF�iuA�����}�2Qڱ�梨��6{�����G씾��O*�I����ޅ���I��?�o��z"����+#���W�o�����<A�ρ�)�U!gQ�ͳE��#�==%X��������Q�"�Μ/�mA=��	�s�i�"�P3@�ݐR}���ѧ���ƀe�?����JF>?ϸ]����q��p	JD>������A��Q�? �N���*�p��|/ۃj�	��v�VJ^fH�" ��׏�gm�Z�?u����I��#�"�qȂ.���t�����#���ܤ2@Bc�[}��~��}u=_	X�]�݈�&IuY�L��&��$�e��q�WT�wy� �.f�]9Ֆp�:�3l��1�U.nG��T��\z�c ����E|'�y���	���� ��@�&�����7�C��#6l	l1W�I^��kR�����z��k�Ҭ�:��M�_&���5j�yvCp}��5t�X�|=��%�j�D�xOW�s�����_�6���A��(�N��@�LZ��p�+N��g�������W��^$S=��D�	NL'+����p]����B�o�o��?��CVuMU�Umy�:�2����V�3=���p+���s��uYT=��)$��C�4�<��:��GgR����z�6����U�kr@���i�w���PyJ���U쥄v���!I�+���v�����U3i$�L�ӂ�	�̟�`�Nf������\u�%NZ�Zi�a�f�=���9i���W m?�������X�"���Ryv����l^�9�G�1��3��%�%&ζ*�>�����3c;Ϣ�ɍ��0(���ݪ�S���"[�����Fz��hmtq��`y��{��*�G�)�j#ԀD��}c/�`��m��;EM�(%jf ���'McZ8=��n͍`d�Dp�Ȉ����T)=������^�ݝS�gh�*Q�6@�mR�Ye)T���i�qP�Eܾ�?�V
��A����$�6���
޿�R�LDLh"�h���L�BR���c���v���zг&6	v�����O{��!�s�
X�I�aZId�"W��5�:�'�Lc��]|""['��O]�!��}��Y�S�Z٘w	�A3��֟��W���ƉY�+������u���q=�����ٕ��u���1JV���>ldF�NP���6|���|h�n�ǈp���)�|&�.����g���颟B�b׌) �|5\w�]m�y�t���$�)J�W	�N3K�� ���R\YJ�@��-���T���ӵ�_�ǒ��M�]ar�Go-�_�L�[DZS�eLe�IWF9C�9��"k�U��s|Q�X�}��wX��(�jb�d��� N�\�k*�i�oo���8����<R�y�E6uY!� k�[� �)xȶ|0d�=)@�(�+��u�4ԜS��2=�a�)KkuDu�%���V��$�i�9�0�#}�ERFQ3�訒R><F�A|d�͸��!�p�� �Su�o����\1r��Y��]�t�1�qKH�����i�A��[\U]/Ho]�=��s�"$Z�\�27�!��`�&�3˫�-�U
�h�ls#+��ɫ��O^ƐwI���zeӅ��#(�<���Q���;a����������P������]?kO�È��g�=�GV�.��7-)^��	�)O�h3SY)�E�Jm��
���g�G]
����Y0���^2��y"�(4����~����hx���`2��d��V�d*߇ny�R�����@��FഺN�hpz4�8�,��P�{1��^�*pi�\C�]c�$_��zNc�����V������\��	JɌq�)�U�	w���u�ءy�&��8CK��/&�BۂJ����{q��K�S��wf@�*�7�P("���(�Q�Z�朾m�Q���_��қ$��Iꐿ�u`�4�_� ���V���.���p�9��4�!r�ok���e�jꤡb���Ai$��M���o6���ډ�b���bm�7^ ��d���Nz��T�Fm��)���"����\����
}���5wv���L��sa���R��IW�e�:�Ц����,����!��v������y�\d*4f���6ry��Dq�k��P���.،�Z�}�N�@ĨR ʅ|������A��C`��W�\Zt���׊��ؓ�V���Fu=�,qh��>p�P:�O�Z�hJ2}�s�>	�<�.8�oC��1	X,�A�&�]�<�ğ��F�>���V�|��G����G�٧����]�T�Bi��g #�?¢��I�ʇ|t�qZp"Dgs(m6��#es��,O�;�dd�������EHsS9��N�v���(��tS�:)��3LX?��lW�x����7�8�Q^MR�*dD�a^%��$3i����Lq�R#�xZ6�Ǥir��eG>�uz�D��;�N�J��[���0�V_�^������u*f�E�w��8EY��oIE�eϝ�,�� �6�e�&),��E����+FS=O�l
϶@B]����M��	���<��!6cm_š��<��l"�L���@
���OT@����AtV$k�w�{8���W�r�������I��R'�ǯ�:�Ar-�[��j��C��[V��c)��DkN��%7n���.Uf'�S�n�a=���Ǿ@���'K�!E����Omb���5�c�x�f3��D���" +�����ʖ{Ab�;��J�$H���|9v)z�V����D�s��,�Əג�u\���2��i٠'�A9����˱�������?�
�zz %�\&9U�z�ƀA\D�Z��ɸ���t
����Z��+ꢬ��7j��M��U��ϱIo�L���M����r�ON�*miW1x���fj����!-:�x�;]�-�Mj4E�i�5�����.���@gaL-��{v/$ [$�2f�BB��bs!�8��"�:?���v���m�Ѥ¦XI'K�1𿊍�jكҲʐ'�r���_ߨ$w�l3��М/��~;j��>���
�2��w�:�F���n
݄��O�#D�<2vED��|4�!6.�z�/�;����U��`�%=�zk�3�����M�
R?�:��w�-�&��V�wi��=�#�޶s��C"�����j�c�G/a�E�z��?���R���x3߹�a�W~�u��`t�AL�@������>�X���[) E[�J%<�6���z��F�j�D������J�KA^�
��Q8���,�)��$�Dj��W�8�`�ؿ�~�l���n��L-6��r��&���
����([7���-ݭΩ'��J>֌�ڸ0D�6�~��i��N�\�3��S�!��%zn��'p�4��A� �c���ك2���e��Eԣ 
6[E3��w�=���;�SOs��u�kK���JQ�L9U��(�'�إ�$�T�9�]�����2M�+�b�����0�<�K՛�Pb��Չ4:f3�2�.��<���q���"�_6��F��o����v2�ThZ��kT��lKc�w��ے�ڗ�����Y*�������4�c�;��3�蒘]b��{~�F��<n=����$�ʚ�ep�h`qy��&�/>P4��NŊaV*{֐o�{ӆo ���\���.r�)�9`��?��h�r�`���R�p��~#����%�����~7_	dC�b�t,:Y��RP]��� c�Vkh|�Б�y���Au�+vRVV^s��eF�߉�!�V��}��7ëog��K�9�-����쿺���-8XHw�Z@Ƌ4j����ܜ�l�`�{���t��x�6�`E~e�3��U�qj��οTCs��S[{��8-�䐯V$�bgu	��#�S�!�c�т���^ ?�1j�ñ�~��oe&� {�>�-�Ņ�Hx~G�!so���Swǵ �E4�����}w���<���{��*T�%Iv�2��p٪��^��s[Oʜ ����&^����R�YQ��B׿��..�QT{BG���R]f�W�Xj�q����#�.rY�e��ޥɿ߳{�h;I��k����Y����`Ѵ�򕕶MJj��`b�MDV�����W���b���5|�{BW"��o������gY�%�a8�,t�����tf���ү�	e*W{Tc�yCt��:K½��u�7D�)�V��B������N�]�� @����
�k>�0�c���G��H�̵��Z�,��ټ+vڨ���Q���ON�6.?���1���M!v�%�V,Ŋ>�ػ
�������5®u�,PK���$l�XQ�&4�����j�^3�H�_#c�m��@��>�t<Ұ�]�9�uw���ud�b����yK�K�:*� �_�E��e� �W3k��l,�f��U�k|�}vu�-n�'���s��N�bx��L�,L(�y���ț��r'پ�l��S�BAU�����k��T%���-\�4<2�H�L>{Ez���4"���le�������y����uaz�:�e�ͦ�\.�1��xi�T�ڛ�b=%aE�1g�w�Uz)@�l����PSʊ�m�ג�v�TB��Y��n,w���G��+�SH�bɎ�^ɖ���R�[�m���\"y�`\an�9���{��,��޵��A'Q\0C��^l�f}IZ��a����.�<-�`:�U�D]��E��J��Ns���4���pk��C�c�K �� ��1��M��������#��TD�R1[�>%h��Jb��_�9/�hJSn���W���fp򂆙_���OZw�z������Â�ER�ŏkz��(K�!���W�ԥ������VX�#b�j�[\
e�ky""6������-�QЉ%ᘓ3ѴR�E�/�c�s��v�R��<V�p�9�95Qk�Hz���=��+)��,Ƅ]�x��z�@�
K7��FH�l�W���hp@�}�M�H`<ҳ�#��p�~s=���-: �Q�@G��C�(�k�5�=T�NHt�����t���@CV�	�>F�x�`�ï����zF >��M���f��w�2���.�>s��8�γj����8�^_�̔_&so��d�W���K7˓�w���&����3�P��> I-M�F�W0+o+A�{���V�4^s�_��ގcq|O4?/��f�@JS|\�ڣ6���1JaFC�[�3q�0M�p��� ���Z:fQ��G�$|��xޢ%(�J����F�mo���ɭe�9�3.q��7�"Xj�E:��������
p��=%(�=�:���Ujz��0d�k��wu i�nv��:�bbi7^���B��"�X�ب��q�\=��=� ثk� !g5��GHI# �q��'�����-��dU	��ʙ������GQ@����~�U�V�5��O�� l^.�+y,b��z�ز�O�b��^ɽ�.)��J�f�e�ߣ� |05t�$��� ��|cyk���l�E�DS��l�L ���R����%(K[�����������3��W2g��J�$����;8�+���B�
xCË��|��d"S�P=I�r��S7F��U��՟�/&lu[Y
E�FT�Z����9D�g�0O{b�)������to:d��.��'�5�.\J�����y�%�49d���Ud(:��m��!�j�~�S+�wd��)5-��	#�J{����	�pwq��}
C2�Jt0(	�o$�
�^ZU�`^�{��lZk8#`�}�&+s�@�+9�x�)���&�U{�9>��ƛ�8Ӈ�w��/���5��,���\/B������z�F��OR*BB# ��-������
�;燹[�n��ͫ�K�,O̊^���Q�~�^+���s��3V�Y���?pi��(�T鸬 �P��A�j�,���W��s_�yB,��p����T[�x)�'��Y��	i���QQ����^],��Z�PVF�EgJ{l�p�"-�o���=X�ӷQ�8�7<7��`����U�rƢ�gIP��µ��)%@���_�n�eB(�*<j'o8�Ͱ9AU�zC������,
�;��>��!M���t��i�_D��A9��M��=��09bOS�c����/B������}^p��#��/�J\T^R4�����28̅Ծ�'����C���'t8S^�\n�Ĉ��U�H�c=|�i�i�nF�Z	Ú����>Vw�Xxح?���=�� �G�-a�)�ɤ�&#���	�QFm�(KG��=�F�����׹4�s���͙��@mU|���
ʬ�6(ʧ�l3�L@6	j��#�5���$$�5�"�]��y��Y���b^8�m�Cd�[�
��x��}�	D�$����*��~�t��_ԛ���X.U6�O�T�Y�$q�Rןˆ��fa�3n�l�._Oֻ��3_	�C����5��2e�[e�!'w�]HC�q��|sT?}	����W �>|S��M*Btnͤ����HEVUjj��V�?�93��*��E(CI�� �׀�p�z���\oY��nk�]8\G�
=r�o���ә}@���`�qA�d{���<641�,^��}(�Oʎ�w?\�rj���غ0m���y~�� �>͔#�?,R�����ae��o�o�߶�թ/�4���""mR�iU�'�O�)+m,}؍�L�݅��s��Q0��[?�$��u�z����礻�!�#״��q� g�E���Uq�Ƕ�V(>.�l1ż��-?w!ϩ����b��ט��ڳ����@t3Y�,�aB�6� B{3e���}懔���핏����1� �m�hז�6/�:	wy ��mp�����h�����L6�X�#T/�}d����B}�N��7�;���oA�=��Kq-"|N@L����H�9��$1��7�)�T&���1F�+M#f�yY���f�'�A��~���z'J�����j戛9�?F-����b��-�F�4˒i��2�T���RU���e�>M �
<���,��u���
d��'{��q�'��,�?R���HB�k�����N�dCu�	�:��k��GC�KTi"r�D�W�	K��(����oD������_ff�_y���P/^��2��'l|)�GϹH[��5�ֳi�A�eݵM���ȕ��,T��.�y��a,v|n��3u,8�@�5��|>u��0Z ��/�_����U���{4]�^�HYF�L���b��$�C�Wi�(ނ��ʄ��^��K�&���_D��)�i+��A6�,t�k,�4��c���HK~h�SyQ&6l�(	:�{���4��]R:О�C~��6��������U0o��d���yOa=؜�i� � +�*������ꁛpF�Zk��W)Tw�Ey���`�Y�� s�J��v���������P��JK9�zq���V�X',w��>L����u�&+�^�:jje���n����0�	�V�қ+
�m�d�x:}N��$�"T;���
������U�(*&�R��/�'&�{�`e��xĐԞ5!�
���-Z�:���"�������5E9+�`�O�ym������@��1z�5����0k�[Q���hv�<'����4r�[�o]�+�\m�&���&���{S�:I�I��zW TDR�w�qԺ�x��E��mSf�� Q�&�=c���B��o}�N2�dj��丘��77�ե
n�u.�Ҍ�p	�ݪ���:	+�S��Z: �1J����.A�Z� ubݘ	������L���u��$^�p��v�KN���0~F���\\�`{��4��/ƀC�N�ꤘ4"1ӿB(ڱ@ߤ��&����56[�7��B������Ű
Ϋ)*��%Ь���a[Eꬩ�ǜ�2Lu�{�+qHdG:�|B�Rk/�ݛX��yM3�:<�nx{�_�,�<��`^A�^�/%gf���Jb~�?���OMA������ā����V����¡Z����伩o��$G	�v�xV�$��|s�t&�=�W�7�TY U�_�Z]r,� d`��g�d��/-�s��óz
���7w?B�M�ڇۅZT�]	"�G��YD+&9Ɗ�'����y��dn�%7�iY�4w����j%�ԭ�
���F�����{1zˊ��y�9
WjY����]-\�j�pTڃit��d��Û)�Xc�U�l�1J��v���oe��Wu^��i��p�9���j�� �O���
D��{����Cz��%0��-�S�Ɓ�q�Ԭ����㉜l�(�3��䉳�Dk��;�G��j�dW�b�������#>�V4��~�~� #&,��T+V:�
�)#���:;��[����.�j�D���=Y�����t�\n�n`������`�oUU�RK�;w�ê =E.�+�/ߴ�R�O�嬹s#�&N��a�wQ���Cߊ�O#j���*��e��B��b�y�zl�Mo�D�8�7��2�שּׂ�^,�a�_�59Q3��L>�K��$���r�Sr�`b��np�G2/C(Et�s۸ǋ���W.=_U����ðW�u�{��+��x�X+��\Y�I���f�v �~l�K|�" 0��uڼ&��@bB���v��D�T0h7]SK��|�P�Eh��w$]��#��~§|Н������g&��0��ecб��>g�L(
WX�D�HL�Z��MiF17�#�g����� ��w�>�a%��R�޻�\-R�r����GN��vS�;��/q[3Pu�0���I�8,Ozr^� ��@�A�F&PRQ��3~����>�ĝ��4W�u¸4Έ�[�?6 �i��>Ϫ �z]�*s���6
��R~��9J�`WB�ll��p`��tqO=Mw)^�@�B�$�*�o_�xi}��|-���4��e1ޓ�e8L�m�-��R�dNX�	����;��.2��	�����E�KX~�}�꽣�H_&� �7<�ʍ�4M~�G+	����Ee���k�Ǒ@WI���X���:�s8U�
����ϓU�0)=�7Uj��V����0�,��A�(�L�V/V<���`������֥L#dp�!#�������s��i]��}�z�#l�V3tt�����H���OX�Qr�BR[g�F�@�{rZ��L�H38I�js�@�y��rB�n��L�OƆ���Q)�����3u�9S���\C<o��fp�5 ."���S���%��]����G�|䶧G�)=(^z&(�j�h��y�Λ�G/���z��ͽB��ڛ^������7Q:7���k:�U>�������� ����ka�$*���Ph���S�9�@u>֎ݏ��@��|�J�%��a�BBϴ�nY�0ˤV̛�Z��=_(;��϶��qe��ل������Β��~�e���?���p�������ܚ�[��f_>�V��7�k^�z�}S˷u���nofT�J=�������N����yl���GD�SK�V�,�"�S��q-��@%������Z�IU�۟Ֆ.5�Llt�KG���񠢱vA��6F���(��%�Ļ(��Bu��[��A�2)V��L�3�﷝��3�8�(� ��y�1��eb� TǑ1"�WB�	�P�ǐ����E�����<�3K�A������ʢ!����WZ���=؏\�p�6_ʃ�]^�׵ph���� �m�.��ػ�~��x�M�s���Q�./��a:��~-r������X*����w�wt%Q���9�r@}6������x˶b�|�p	{@;��EX��O͙�B���s����@�w�-��5q����`�k�݅ ٤o�<ۿ���I���H-�M��ѕ�m���ei{���"���{�_��7��r�O$�^�����U|A1n�G"@x�4�mҢQA� �u���~�a7�x�R��T�*E_<Opr1w�pL)�<]/,��C��W�8��;��T����bĸ��DO�d�l�Q�#�䌺���pe-W��O�C&EI�CG�F�	�xS��۽'���F��t�m�_?0�1�p�kW~�1)�|��y��~G��4h:�}�aͥhU���v.��x>"��D}|.��v�䘵��? R`�#��3�L����"G�
��P�B!�m0�ɅEG��L���	�˥ҷ��w#�`N*�()Qԉ`�-U����� 6�åђ�Z��w���-�y���*�u������V˕j [',3A�gHMGou���Rm��))��!�����ę�CpN��䑬�S�;�i����)$O��6�~y҅����î`.҃�������GȭJǋr|Xk`H�=���͸�o�\7�"9G�L-�5ʺ�_֠�E��G�E�d9���a��gJ{Jm���Sr�`϶��_OB�
"Uc.��������YN��rկ: ��*ժ��pl��Q�;`J�[�7&��#��� �d(3�������H��-���Z|��N�v��%��R�ӕUu�0#N��v�ApWkL��!`b�)]�2lw��ˋM�K�wݬ���MBO�#�f��I�#��oX��� α��2:!$������"�w�0�ނp�Ng�^=�q����؋�L��}{�6-�B6Z�b��
/U�1���'�f}�; Ѝ�eۨ��w�SW�0Uqϫ�o{��5d�_��+�|�%�����L5�5yz�F!��{IO�y\�����X���I�yq�ґ��n�x_k��BI�0�m}���Dݥ)�C܀�9M�R<+3`��lmd������2{bsT�t���y�&
�	�frՍ�L"
^���"7���i:�5dӊ(0�����n
��7>r0���5p�bc���UYS�7�,و���'Pč8x�Q3�Z�h�obt�?"�����!�:��x���fd���?|���!�,��y#���r|U�h�/�9�zà1���]W�~����f������k�l�w��/Pez;�r['}��p�R����M��-y��nt��U$��I���6�ʠj�DRΜ�Z���ez���h"��z�i-�6(GoE�;�% �?ew� ;�|ʔU��/WO��T�z�� j%K�����n&4j�E�yo�bߢ�d+����W��Q���nW�whR`L��1W���Ŷ2���OD}rW]S�ʖ	�0+�C��!�Z�mr����ݎN	.E��'�]����U&*�>�sQt�e)K5����	�-_ ��nQƸ����y�B�Ao:u��]=0�����X�D�ݖ��s�eU�M�_doﱩ���۪P��1�����۬���kf����mq�@��'�QuF�]DJ5�I^��7�s���EӚ}���Z6ر1 ԩ~�L��쵠21�������R&��
gY�u=�ӵ�kU]�^�Ǆ��b�
�8M*7H#�輻T�v,/ �5�EF�Op�zN䁫�ϗ�t�6B*��9�+X�2���T��x��H��D���D�kJ�p]r՚�xyz�.���G���{����ʍ��o�
a�>������/�'g��6?JW��{C�nC(������z�׽Uu�Y�`7tG����^���,.A&���z6B����΂���ET<K�v��>��I��i|��D�BJE�x�6c�.Dl�k�r���X~�>$����E�
T�硵���=���C�~�}Ql`Ԉ,��̥0�|�2�(���sK0K4��ƞ��iw�itx�T≾����	^�j�q�����t��ݒ<�Vn��4
zԥ�Q�����_[��AF��/�S��n�x�+g�a���f5�&�K,�-�^Ë��
��~�Ґ�� ���bGטk�@�['t����wYX�'�+f�~��P��Ľ�9�Ua�%���Cv�������ͭ��,W<lB�ĸ+#� �� m���҆�/�E�`�9��C�*� 
N�����5�	ba쨛J�uF&�$_X�:�	:�_�$��/z�`��}��]OewU��L�޵xM�X�]��6�
R�ԲR�~N�fK�!������:��-�5v�����X�������b_�t|f��֞ �tLA*U�ys!T��کyn�ۍIB�`�m���3�=���$L���f���n�k�o�C��N�X���[�>5��C���g�8��0������:�/�@0���y��&�$�F��O��2�_,.����N�߻T��J���A�M�NO�ŉv��e�/6"�QQr	�1�vBs_��p��L��\b0{gFM�3�$��т��a�����P �F�5�Eh3S�ص �8�Q��]�'hs��}{0sv�;�>΢7�­�T�����NhIk��g���X�$�b0�8�X��M�D��I����y �Z.,::��O�(��=�'A���
L�u�Q��	$��C��o��Gg�[$2��m���T�N�hB}=��ܐ�w���w�����2�`Kh�}�eZ��J�.���1�������]�T�b�]�l�p7�2�N��dX_Ǭa���o�ѭ�|���,���8���8��Z��=T=>���e���i-݇�Ѿ��\u����:�!��H�b_ԯb����p53n����<QR�%�DQbK0R�M���H�p񈔆�[L�M`�Z�iD�Sj{�c�{�S5D捺'�=�B����Y��[���=E,	��=�/&se�YL?��"WZU-ҥ%��?��M���8�����	��5/�k�;;&��(A}ED�ґ'3�r��EZ,ύ�(��nCW���$�Gv�V���O��P���Ev~P��l�l1������7��K��&i�;�!X���A�3�%�8�F�K^��F�a_pb��<I󍫒�x`8�#��PQb�yj0TL��z�:I9��!6�q�y��
`�H�<C�F8�=�B��K��T&�o?oz%���T�cA&  ��T��l@	�����^M�%��+0�n셁��dh ����M���<�M��9���j��]GIG�Txt덼g��=W��'���Vh�M�vX�Vf ����f�I}����w�0��Y�K��6�{�۸t0%�������^�Ձ���л�L6s+jHG����/�z��eF����������w9�[��8%�N1�V�J��;fj+��E���`�;���Ґ�h�៙Hi���I���^p�������a5-���#1��P�N�/��X�}����x�Y��&��s��A5U)!��ِh�޴��?~9�&��U�b�ھ�~e>�)C<����)䰯2��&&&9������ja�~������߀��t���a>�;T�u���;�-�����%a��//�Y�xʠ�����,V��V�*�[�#"����6����'cg-X�\�3�{C�qs�����tŊ�4��*�o�L/ԭ��Es���R}�$�9��ES%v�qp�C�\����Y�y(��65��\L&�M؆(>2F)�R/�7����x�dn?H-)�;�P�y���%��T��p����:.��Eq?a��Q�;1.�כ[~8�K���{����Ԏ��R,�p�x�'��o�n)��_�~q�	�,���)�*�����o9��(�&,z���܊pQW�@��b�>�n=�����]-f���@�H��� t�O�~F�̘֑"��iA<�}��ą���%U�⸊j�wڛA����ŧ_ɸo����0��y����=KK4�S���p~/z�G�7�p��!&��/~��w.x"�b�����b��HFǡ���x��@�aM���b�aTt��bL,j&��e�dLw}�.+�5xGŦC�\'�:�Jm��R�I5���OW������M0�M����P���ؼ����`���SdQ�2C��d��j`���gR�
el9ץ����RpsT�\�[���J������T֟���x #�n�h%ĺ`UL�'%��Q72c���t��U�Ba�@C����>�2ԯ7�
ܹ�vꭲ[5H�:j�([D��[]n"y�!Q-695QFf�-T�q����V�ޟ���Yb��Oe6���0O
Jڸ��rf�P���6�=]�ЋK��$i���:KB>��y�N5{mItEK�o��>�7	�҇C'b V����1k�7�I7�X����I�P��.m�@���_�p�$�a�p�F�G(j��n��)\�o��e�=X�%��P)o�����G�J�5I�S:�����=�S���F�9O�{��\%��7!�:� �����d�N��G�a_�0'��\/I��:@��0��k��ω�x�z
`Fa�]D?|6k��i�yH��J�n�(ÐlR��[1�A�E7$��꼝H<_�Z�z�
�%QV�IASgi����뗝���b�8���7p�LyQ
2rt(m�>j͂��c#+o��_��G_�5<	��"�uԝ�5MY%�:�ܜBcn���W�QM�Q�����#�����T7���V��RvQ�o��)qd7W[�{EH�Ѐ�ƛ�e+A]Z!3�_W���[n(�=�]�o�H:��?�%ķF�
B'��W��k���BAU�~N�k}?����C�g�qy�k��ض��Q. |T��c�<:\ا�
|a�/T�z�3�cNw6�4&������``)�]{Bg�{b(y�?��Na�w�2:9���ot�	��pK��͖�B��-M�Қݥ��=�m�"�	 ��}��4��5e��m���aM��ZvM[ݗpP~�����a[�K����{�;�Ά#��K�}6�xq�5�ޣhؙ!؃?'�����-��ы f�j�~b�W�``#�=wOe�����Avc�B���(*��F�bq� ����[b,�<�Q�8 ��b8PC��#uC�	���3�5>�I���\G�.P6�[�؝]����6�n1bj|�אk�#1��[La9��[�]�v��#�W�az��XÐ)Ho1x GSȔ�r���~Xs��)yZ#��&V��iI=(~�ų�c�%���}�,�|:æj�t�GEehߪ�D��׏/�Џ ~�#�w0��.�:\�&���5�b^����P�����;������
�)u�.�S �oQ�7ǛM+؛���L"� �o��#���`� �^y���2�9((���"��(`c&����
\����(o&~gO\h>ٷ��c����'=[�?B�&��s�56�[��p�X}����D?7�SF�8�idƛ ��\q�i�R��3�W LP��J\�Y�LW&ޞ9�#M�c�q}�7Z =A�4�	�m�U����A�o�@-����q��~S\"s�&օϻV��`�BZV�
�"[�y��+��FB>���1�i��1\S�3d�_JA�����+�Ҙ�u¬�)�D��m��q^���X=)��o4��r�
E#���7����$d\�6��K�s��J���Jp|��܋�>�@R̞!�#�K��E\�� H�d�@�`��B 8�G��{��2,#�Ε���o���[ҵ	��!�
6��[x�[d��zv����9ϭۀ� d/�pȷ3��EQ��}6e�`��pŝ�6�7W� �����X��b:�t�Y��xG�i�1�*d]���kNlė�j[��G!<�#I�J��[l]WS�Y��Y�{����/�]I��]�D�p����R�OC����� Ǖ4~�MG����1@��D*�
Q��C��M����CU�ƫ��ٱ�*]@l�Hy�PK�]���3!;�8��1{�7����x�J�H<�˼�wD#��b�I�t	Ǝ���="��1�r_�r�`mk�8y�YKo<b�o,H�%���ӹSԗ��l�}E[���z��	��AW�X�E'Έ��ЄGQ�**'��'r���"�����fDX��M3�1�s*yS'e���J��WC���s��]�n.�9{9�7�h|�H׃���5a�L�?&&~5�@z�����m��o��9��U˾��i"i"l���}�R�TH�p��MB�} �s0���z�$6�N�R���-CKJ���5D��ׄ��#��`k���x\B�|k�D�Οz��i�5��j��T�gVO;o�|�@[ň\ Y0�LOM�����C%����"4�Ŏ�����y�߀�"��|�����������K����(؜6�e�)tλ�;
|ԕ?V#N#��K�:��!�˞b�
�j���SL�k�d�P g$߻Jof>x=u��I��(���7W'��eo�N,k]�C�2��!(!��Q�r�/[���<��xs9���y{Ĳ՜w,�rBb̿k�@>��ş���S�_F�Ba��.9�)լ��Û3����I��>��'�#W��x���6R~�PS�kI�����q�W2N��}����N 8ރ���m�������Ĭ(��	T ��a���M���<u <�}�O0;�|�}[�zI��n��!(;�����o���A&)F�&}
*y}n�33�L�{�pe��@=(��[�W]]ڙ�<g�r�#JV��2����A����I�jlf�*�OTYE��Ay[�c�µ���l}��a��X_�9�DE ��B�h-(�5���]I���ڑ����P�9X�
x�:���2OE���D�LC�WkK����i]D�3�:�|x`��Osl�o�<V�����X������oWnj�����Z8�Z/3R2�i�G�V
�GJ,�M�7�E^\Mդ��{8�%+��U0�a��&��P��+����(���n`��\���We��ѕ�t�4�}p�DOK�R��/p�cX��.:㦀;��Q�G�Rb��4"5HR�I��Q�SG�5
l���L��媜�Y�� �*D��"��G��\���u�����o\�o�d�KΖ�؄��V�Us��X������V��oE̛o���d�7���T�h�A7*�Ј'�tk_��+��>����^:*���b���~oW����%���7;�g/�i��"r��&B}�iۡ�>�(5��5�&�;~�Z�������<fͻ�
,l��?$���Sb�ѯ�c����9ֲ���3z<-D���ԇ��3��?�e��O��)O_���2|6�׶8���hW	|��F/�q:�U%&��/d1�(�s����)���*e���#2� �q�`���u�T��`ԉAG��-��eWh$�!���F���E�U둧"*�.���>�E� qjC+�q}[���H^��f(;G+��x�n}v� `9������&��C7��5�2>���o�ow�X���%��ND_3am��.{4�v�����z[u���ge��		�>�\����E�!��r��b9F���$�@hH�pN��2Mᰅ�g̃x2x �o�k%��B��KRVc��������f�����4wl��,��m#M@M��J8c�~��NΨ7Xbg�~R>i�VA2�F�[2�ۊ9��T0'9D����{����r��K�O��Ee$\����.KU��
����ٗ��+�_t�y�&܅�*�6����F�xU��������'�E�1�g�%�k�ʶ$�{�x�O�%��V�U���Y���W�_(w��G�/~+�'-%#�~u2�k��a���5����y�^@ӆ�ʁ�_6ɂbQ��i��E��z�S����5�R���\�3�`z���g�Q?�iB?"1��+y�{خ��6��0[b. %�����6-��u^tKW�G��f.��Lߘ��O��a=;��8S�	�G�`T �?P�m�0h�- �����*$]�9����d�g^f��1�z���@��O(��R�(N1�Q�r��SҟL_>l�7�W����C�(Nj��~�~��@�{t�+l����<��P��)���ר�*2c8'�aݑ&�`Yy?�xO+��]��Kf�碗x�@:v+{�gO��Uէ�@!�t�Z��Z)��3�%f����_�P��vc4���.���>ۧ*SjUa�w��X�L�b�<�&��/�Tԛ����Ų:��3�o��O3�Q��m���侁K�#�������g$���'����	��J�ꆣ"�p_ ��� ��7s�	W����D�EV�ΎY�Ǒ�{Ŀ�b�?V������X��|&�l j׬��y�="4�᫋�����V�����cѢM��w~�l:�C1L(($��O:~�M�݈$],�J�	�:ڃ��G�o��k,ޟ1���@�L�tk��U����<yk�ƺ��"Bxg�`��]�Ymv���[���#���!�x��J�yWHΆS_�B���]�D�������t�}�M@ ���d�Yͥ�I�C �O�0��eޭ_Ϟn8�?l��h��5��H�����˽s�����1k5�@{�VF)��k�?;l`��o1�<�>TBw��(�:5
��b�e��r�ުu�C�Yo`�q�ÍW�e���c�\ƨOXrZ~#昩ꏗh�ޏ��_Vr�W .̪_z���֌%+{L*���Z�H�*�?�n���Ek��3It"�������C0Z��i�E�>���NŜ܇0s�esA���8(�����G�w_��0 	i�JC�@�&���u�#�G{�$�'4�yk�<�'��V#NυX�p��د��Zۘ��Bˏ"�KyeŕC���hn�(�1�����!��+��=�p8��4����_$��v������I9v�l��"
����?�m3h�#"��N]"�39!w���w�L�I��=8���X����PAD���J��
=�/?-l�9B�|��u�K�Eٚ��Ė�q�����!��͝�M\�J'��aJ��g���!�b_PZ��q��֞������$�"AA�ED�ġ�A��y�*�-�cr#�M�����h�o�f+�q�=����&��n@+n�Z��}^6���ga�Z?x\�a�k9���c,�-�1,Z��5�6�d�>"j}be���.�zA`b�HH�k'�k&a)=��+\���"O\s�#Bq�Sz<�"����9ZM�;B{ǔ9s�	c�޼o�����+AN��é2� |�9���"��u�����9��
#�]ά��?��7[H��R���i)�Ӹ���ikV���X�
8��!c�rN[�����c�ab�C��8��v-j]{lpH����\��jK]��p�H��0�J[E��������FR&3�O��%���ݕ��:q�kF(B,�G���Q��b����u��+H�r�G�aaj�-� n�W��k�Ӆ> C@���eF5F[_&%�,_�\v�0(%���<w�l�����CQK���CM΁�w�M�&-�d�PZS8o,��͡��Y�-�Q�;Fwk9�}Ɍ�1�++���*J|�/"b�!4�5ְ���& 5	���ȋ{��H��L5jkj�ʨ�C|�i4zɣ�|Su�����Q������W�C �"�o�n�Dw�~�iY��`]k��ɡ��7�ڝH3k��'��Q=�G�kEunǘ9�pO8�!.O)7���{aҞf��sI\-�sLED��]sʍ���T��|.
Mf
���{pí2n�3�ν\��:$4��9#�C�F��4JI�w�z)�L����=��S�c�=l^0��]#0�������"�Y�RC�߈o�W��^��N��.�!��u\C^���	�@�
�eqnw.��Z����`JOB���D�t)K������v,J��ǥ�x8\��q�-�`�>t\P��G�s[d斟R;
=��?@�2Y.q�F��6�Z��,k5����V��8W`����!6�:��)5�.��B /��x5$v�"�V C]n 7��(�VTR�f��Q�D~�[q���|���)����dGAU��'V����f������Ο�,�Ӧ4z����8e�;�����V�k�<��vXYH���'8�n�� *����Y���~��G���͍�[�18t��t "���VAǱ}����Q������Z�NA�d�	*Sީ2�p��eZ���~4�sQ�SIh=�FN�*�j~����.�N&i�\1�q?J�,���}�Ap��g!���߳ud�
�?���d�	�fR���?.1�������O��	#�7�j��4�\#�S�t���M������K��#��9
�+�������Ы�)n1	^���+e��Qf����,je�Z&}�%m8�&��{t*��e�Tt�δ4��N$3T��r��4gVI(݆$(yI�-Lg�R`�w�s1�r{\�fK�7 {�F4Š��ǧ.T*���|�3���q���aEun«���W2�J\����9(��d�*����&�T����������:n�G�&q�
v��$��a.������Z��b7-�g{�5c�?��C7�Z���ژ�+�J'��L�w�Z ����
I����~(�L���5�m1��ۺKK�����T�@�| �{5f'�<l6x�d��lH�侏D~�,�j��$Z�u�7�:��5X�Y����紇.O�:�b��qm���.�U|�:�T=	�D� s3֟Y;I}��m�Uٸ��LRvq�M��Lc�X�B�q�&��6���|��\��v��V��Nx�*��G-�u�<�ʢB���*$�#wCY�Ȁ2O�i�=�?�Fb#|��j�˳N��gR|ݪ S�l��lU�r��ԍ:=�{�����%�!W���)�kGG�!����h�Ԃf��������i['C���pwi�'�v�<��0a	L�o=����6}�sU���*D�#�DWِxzE4lu��H��Ym�����@�t���ň��\{2@�ߓ+�z�=�Ù�$���w ��s�*GT����8���F��a�J�B�wkξ�5��]�D����D=͇�aᄴ���Uy������Sy(b��`�&��3�мJcD��p��U�![o�L"�f ʁKv;vޒ�#��������n�䁼��}Lg��j܀��s�hJ\�ai���Y&��IA����"�|>�
au| ��9�	�����3�x��d"	����쀙��r*��,�(l�Z�!�P4�,��er�Fkc�L�dU�Q �F�jf2!Q��6�7�tWs��\;Ŕp�E@�����եn�7"̞;s���w�~G�c�]X�/� �*�˗ȼ�[f�Y���[��V��i4��j���	9#]���+��\ц
q��4����*��<��V[�ݬM/.��%޽}K�AubxD791nL7(�+�;��<�I��	y<�5T�	�cC�(��g�4���vOL'��I~�H��
��0�~���]���<��ԃ�!��u���ZMTӻ���"���_��/�/&�+�l�l\ ��ش�ˈ�zO�Oث>ǁ��]���e�G�9�Ϗ��S���J�F�>�`����α�Y��~<�\S�o*+f� ]X���Fs��Dz5��O_[�l{qu�BQ��.[��{%�j���F�8��|���+�1�JM�fM�'Z;e�:��*�����
�`�����*Q�
�<��W��`N�
��4/do�= N��K6TV�RAy��B�S��Ɯ���n�)��-�Ų<��>��(K#�!-2�X��-P�P�f�������ԏ)&l��P1�����BY2��s�v��.LG�"{��e����X�B�H��(ŉ��u o�wƄ�k,��U��1H���[�?��*�����a*�ܠ8iHY?$-�z�ƻ|�8 #C�.1��yN��D�у�J"���žx��P�-�FXb�\K2s�=� ��T'/@9Z��ں����������J��[�'��|��RL�q6P6w����| `���iT�N5�?��'�ց�������5�'�մSI�2�JN�#{��=B�0Px�I�xĮ,�<�e��Gû����J��F��X��	���������}���a�[T:������.^(��b�}�t��*.{���|[�åg��^����G�"����j
�`�|P��E����`���VT%ۣ(�XD��#q��t���ݨ|{���ώ��� i$�_pzA��Uڸ3��?�����
�!�F��g�_���������>���~\��ӏ�l����6��jؔ�ƪlЍ�E�Q���b՗���x2����P�8�vЗ��U����(�$n���o�Dɰ������B��-�Vz�a|���k6|�Ы�ڂ�t�>Kby�삼A�p���Tx��%P��F���6�%U�P��{ٜ��2��	v��$��A}Υ�C:˵���:�7k���-c�[!�s���@W����[a�>N8��ZnH��ˏ!nl�?ɢ����\�n�J�X?\|��;{�c|�����]F�E2�῿'��.���ZL���TjY�꾵�Z��Q�)Y�� �W>�Z�c8b���pI����6����a��ϬZ.���^5д���YF�eǠG�e��(��Jc� �����L�-��JWڮ�T�Y���:�	VckKP*|�;,4�����������<�6/H��oU�I�T��.n��q��(���J�/,��CZq�Ô�D���f��������>�J�o��`Q��/YړV���a��x�PL�E�������4K����DBDSP_��B�&����&�P?��N�=0�+��4�Dyh����o��9	
)�pdz�w�w�[W���_M�y>;K�H�c�\	��M~��L?�+�K��A���(�r��Y\%�:�q�M�{�G���qݐ��t^�\mLR?�QN�@m4�8�p>5��>�"��?4ǫ��<ɭ�I�k����w��;�>#�Q�c��v�4�~��ge���}���3r��T�A��-_���[^L��F��x��7m����p�-�L�v�)¹X"��?L�����3̐�dEH<��Y��i�X�w`=��L`��+�q������3}���~5G������>V��s���v�Uٗ�4���+`���S<��=����|Ơ�9�]c���$u���ۚȜ?�D1TSA��%���M~����@;2�s��O�$�.~F]���K;�|��Ð�H��$#-����;�J�"׻��ҼM\F!Qy�ō��3yW�aYz�M ����ȑ>_+�S�PZ��^V�.��s�����t�UqjKg.��N ����tM�]���Ve��eۅ12�������y��Q3�bs���(M��f~Y@���l�VloJ�Z�M��n#���ֺ��2�IDp������� [XQj��51�6����Gy3���=W��7ί��"��;
�jd���0W�Я�t*R9�~����X�%I
�2s�r�@5/������-������Bi�Y��S$��:��bz����B��͎๘E��ŕ�2=���)[�!O�S"ŧ�I���m]����X	b~�j��F>�GQ����Mi^���Y�go!���Q�z�R���gt8�y���7S(��"i��{s��^�3*��������Kƙ5�Ն�R�κ�M�XSIɄ�d�y���yO~?��#w�fiL��D�7B��KS� ���)yq+�lk|�r��W��T#4[�15>���07�]2C��H.����]�k*��*r&��4��|�H�o��nP�+S�@ @3~� :���ѐ��<�����,�6{�%���VG���I��[�D�<ZC�eHp��ܭ�e}� '�遈�_�s{�6��wu�T
� ®��BP�c�}��O�Աc'Ѵ�ы=�ޛu�U�Y��$��qҊ�jτLmFJrփGC�~gQ��;���]�G�o2k��X޼���pv@x�`
d��"�P>2�q��鲆�w�� ��L��W������x�0W�缫fa9��Ik���Uk��^%�~U���dT=��H�7��?� ����0%?U�����h��i�cڣ
��C?7 �|UZRH�1��՗\l4��[����������f��"�^9 4����*¢�A���^���};T���J]���D���	̗���<�q������h�O9�7�RKd�zh.������|^:��px����X�U��kXV���AN��h��Q� /�D�X>u��3s^N(��� �F��g��4]+ͬ�q+��QR3�����0�c��
��=�K����V�� �/	ߴ���>�R��7R����3�i`,�V�7V"�-஋"/����HJ�cɕ�_7� nq�S�Yje6�#��h�ԝ:lo5�%�S޾5�����.!�~D���4s*�"k�.�]@�4��B;zu_�L����{ �w`JQ#N�{r�Jsb@G��|�qWN�&�����Xni&*����ߋ9k꿤�S@��@��0�x��%��6�F� %�&)Y�9�� �3pé��f�I׸,�,���-�u�V~,�(F�vA,Wߜ�C7��{b�2eb-iĮ8� �g��6/5:B������=��$�W��sS���{2���1�ڵǆF��Y���[�Sr G%kb���fٝ[� Bڲ�:]�R��y�$�?Cd����DB��s��P�[G}.��#;"�Qo��]y�).o���_��{p_
6�N��Y���c'M�G�;��_ϸ���\��P�E��T���]�G�,s��,�^�:?�K�,�k8��޽~�&o�+�3�6�ǻ#�RC��0��Ɥ����~<"lٔ7Y��]����#G_�@P��\"����)Wy:=|�W��u#�Դؤ8�Vf�[�b�v�4K�}%���9s��Ho����EET�<���{��E���a��P�)����_��j��Fe�4ۨj.u}p�����].��,
��8H�¤ #�F��m��6�Q��:T���k	K#�&|�A;GA5���CV1�a��B�"���6�ѫ�GH���ՙŔ�~&Dn(�DIӘ*�〪�ß�VFI�8�͟鐈��6�ݖv1֒�aI�^@}6o�]v҇N���c���{Yf8���l����֎�@l�Ъ��`X��Mx��\~
ɳQ5��<M���
7�[���J�44�ne�~��\;���o�q�&*(��͊�F�to��+1�G�+}WD�G4��Q<%X�SKH x�Sӻ�&�5�ّ�[�p��׳�h��P`�R�t�!�	0|�E�R�5A�$_Qlvw{�Q����3�z�$咮uw�wb85Y���We�9(�ظ/�$d&5C�+�� A(=T�Z��}��շ.�V6�o:���.dH�+z[�^ۚ�:&�R�yT鯁9�b��2iQ_��-V9���Aq!fr ���ۅ�8�f���E�m��w�z�x66J]�B�#�
��Ǐ�����m��~q�3�tn԰�{�k�-*���Ӂ�U.%���Y]RO�k�����������
�qU��ڤ�#p��g����{��US�<���8��<n�<��Xֱm1�� �n�!ۊ���]��}�l�+�☒XA�-$��ƞL�qħme�bH��jEG�鯽���M%P�w���B��h�2=�֨� P��u�LCuS]ĸ������-9�u"[ОsA��UQ�I�8s��q.b�7��V�ӣC� �������2������z8x
���������j�m �߫G��74Ճ��~Y�)SIZ��Y˚(R��� ��bl�2��%q�RaA�}��ګ F�t�4�u�^��'��N�3 ��<�C�M)+�g�n3 �n�������n�T�+>��f����*���!&w��������_U1����	����/�����޴��%b�xW#�m�fÔ.�q$譁uI1��`/�=�<����}t�8��qI�� �-jV�;�D}j��D�j�K����x��*3�)� ��mL��;fW���ӭ�+�ҁ�2 ���(� ut�e�$��MGzͪ���i�����a��?0�_+�Z&��6���(ګ{�͔�,ׯ9���j)�f�1ls����l"(�z*�n��u�|��sg# D�Ψ�W�'Y�c�P��v6ۍŴ}�p�\���*YMUgk�0˾S��z�6�����s1��� )M�rh2�y~0c�*n'E}u#SF`g���n�a�ԍ�]�����T%��Յ�����?1�Gݫ�;��J�c������Jm9X����xT�d^����6����� �zJ+F���#����h�\�T�4 �)�	֙��O洖�u`w������ۮ�mg��l�9zxH���I$@'-nq�@��-)cw�lZ� ��4�F�+�İV+���Y�דe��C��e�[8���<ؼ�|��O���A�߉���^�|��T�b*X�4HA��zp8ຢ�U3@��O|����^n�k��(S
hI�'���1����F�8��		�)1��ĸ�O�Az��	�cTЦ]�}��Ys~\M�H^$t��K-�uN�H!Ԟ�P�p���{���!�o$��l�	�u�六i7���{D7ド-���^��QH��"�FL�����i�.�ǼFA}tY��v����6��C���"B��ح�*^Ty���?{�2 �>�@)�)�*g,�`������b�����x�p%k�`U��w�2oS�^�d�q�����H�/�*�%��F��\�TÁ��fn���u�YwtN�,�q����-f�L���BaS����wckc��h�?%o��A�,<��)�N�U	5�*T��?�w|�r�/�}i�8�Γ
8K����?��'е�?��!��{�݉�b�V�%x_����w��a�E>�T��Iv�6�f�nh@.�@B��K�_+f���/ߟm2�"�i	�"�I
�O��ڋ�Ŗ�0�=�4���� t��,�J���U�� R�0���>v�ڑ�@֔SC��iG1�֌D�ɏt@�(v��`D�� �ʈ��̊uq�c��f��/��'Y�w[��& G�C9��䰶��rp�\ݼO��9�=��A�Z#��b�f+� 4|	�*���t�&$0�pW�L7�����7��C!er�I*���Jb6���_�x��1��E���w����ʭ�!=�.�V`�� m�M|%O���A8B.I�`���c�#��m+Y� �E-��jj���	���6QXb��5+Ұ��|�kk�&9�7oq�0߀���b�Ɋҙ�?*xò���9x���g�� ����>e�T��e�����F ����|Q�o�U|?ܝQ� ���)@����玓�:���k��$P��d�l2b��0��g���h8��9�h�y5�Y��rBR9^�B���HC��o�㹶-=��a��ua����~�ih��
Y�5��b��RĄ�㍳��tHH�i7�}I�qG�E?�6��]�� �jZ֟�g�`���L�w�5 F-Ϧ�L���͢n��Ar9ȋ4����)X��-�v�����쌫0���A[��f���KG_`�9@+Y܈�ȋ�Ź�aPN����0s��W��\fsa�pq0kW�0�|Kfd穀"�Y��)�)��_M����Ӑ���š��>Mh>`�:��Ҭq�=2�1I�<�Ɗ�¦���ɳ��P��s��C�*��B*��������4�H�GJy�����p�Ҫ���?�n�(�6���/��f|6��:���Ͱ����#y��
jA{"�-��aEk$�p}��v~-d�)�92�jAvOX�	�l��lU
��9*y�KT~c�qa��P[��>�/�ۄT��}pa^����g�W������$��6�$�\�X����5C�@�+c�~8�D6̮_n| �}j�_�˟�L�_Ɩ��>�Eֈ�/�t��%(�m��ah�fR�n$y���&�9zA��[sװ��ZE����V9ǭ�䨃X���Yqm �Z�h�44i�=�̴�-O4g�6��|�`L���T�,�k#��%I����շx5΅�����7���<���Z�������ې�q �H�9�J[�:���GG5�F�v|�M'��jG�/��X�l�AkZ}�l���2�%��)e��X��?��$������ц����y���9�����
m#m*�:���<n3��^�c87�����+���#^�Օ�Ҁ^R��>e�%���{|�U(|3�\W��<Ϯ`�Ee�V�;�=��>���G�Ͻ!�(�L�S���ؾ8���Q.�GK����x"	eZ*�wS��g�P"�~�R¨Z�_��bq9����(��<����#H�@ϡ1� �4O��jp����ȤT]�^I����O:q�U�uY�ӛ�ʁ� �՟~#É�`�iF���1EE�!����u���qM?�e8(<�5�Q#��+���xU'�t�̘�-�ڜ��c�œ'e���N�X��'߷n+�k���o��)e�m�P(����5����Ӧ%,-�i�����6�%9�5�l"y4b�;Sr\��d�����,&�]|�HՔ��d��Il1���|s�cu'�F����[�%xk|�jcX��Ѭ�tZ X��y�2ׅn8}S�ʗO�&z�����F��*��f�Y���B�X88;ק��oV!V�H��x�_�9��f�[��X~DQG�>5wϰϣ�ր�!�$d��B�ܖ��Ţ%�^m���m��ǜ����4����#��X(���o�aД�@S����t�9��a���� 'UۂL�!�.Wi��1����c˺��@/���]��_�6ұm^�f#���1��J ���y��{y�ۈ�!2E��̓�L���w��z}�s{���U�H7�L*~����-���"7IH��� ��ł���2Ԇ_�F��@����Yu�=�'{�v4�s={���5�&�E�Ӊ��~;��϶ݐ�à�;���L�G��7�5?��U\Q9XMtJ[V&H�h�6��f�z̾6jW�9�����F��[ƺ�����桄�G�}��b��W����N�m�L�Dg�[z���'����,�$��MN��z�����.��2y�>+�r�v�n_�o �%��/��Gva,�K���SӕD�G}��-�ha��G�UX*;"&��]��Q��f����.��0P�Е8��05K�y�Xn�h��D�����	U
�~��"7][Rp�k)�����%-� j0'�r\غV���������|�xu���3;�P�5'u|b`���� �	�������Z�R�HA�����5�sh0�T˻-������<�R��[���;�B��b�%�����)͐X[���6ȿd�F����(ع1_�jBC��W�� ��� ~���wA�:�c�6��	H��t����Q=��H�G�V/��8������"(�ͨ���r���]`H�n��� $�?=�HAi�ŐH�k�m�ɖ+�W�z�P����|$n����Z;�1��+��`2ã�D��.?]���E�K�g}	�
����8%fB��:_�P���.&v�/��Ljn��� ���YT��E8Z�~�&��qy�ߠ�
�k1��/�:�� I�{��f�{��#���[��X�KU�ߌ�FN��c���'�R��ښ>�`�t�ì�`K�-��]�?�*|���!;�8%�f��Ҹ%�Z�g�7�t;��{x��v]����o̤g����z�|�;��۶y&M-� ���� /��SF_+���O�+��2�W#��hZe�{�w�ꝛte�6�N��˧�(�k�mJ3��Њ���;�L�J�d���A�E�x�N$��Xx#��q�qn��[�C��hhe̲�n�%�N~S��F�?u���Q���������� +�	6Eȝ��.cp5��͒]Q��"�T���GbX�l�s:���$x�NP�Lń	V�.oӳ����U���|XBn�
M�� �x,�3��;J:���(��)1�O^I�{?�e1��>r�ta5G����F<\~O<�I�hg?����?��%B��<km��U�VZ����*����V���[��P���H�ΰ����-���|F9����ܵ���O�ϔ[)����'ӭ������8N)�QD�V|3�����},��f�oE���OD������k]��['��E�5m��)|����ڼk�����e�Q�I���(�~D�/�����\�>�oWFg�X�eQ�'<���S_���*����ڣ;RƟ�ͩO^5����;��fV@��	�������DN�e�ͭ�K��N��q+pķ�\�j�4'�I�ˊ�Qs��[N��KO1 �W�"�7p2�LG�D�x��y7�K���X֩P��x���I2���p'&M,ؿқ��m,ӵ돞1#�׌�\S�3�<VOԲ#��!�(f����d2ޛ9�/�,��^ �&æ ݈�v���2�nA���on�A�[u�����O������#(��*Qn��~B	���O�[m�d�{�+\d��?��"Ћ���ЩO�AB��{^1�Y�a�����f�;�!�۬ �)ȳ��H��G�r�t5x�]�`��ub诖�A֋��_�[�Ŋb�EW}�Ԏ��㘥� v�~����QқӴ(�To2W���Ⱥ�&��-�Q�7���d������
����UTg��.\��DØzt���5L�1������]P=`H�L���K۾�(zɀH�wi��`��B��������@v�W�������j���V���UMA�̅6����aꕟ����Y�Pn
 k+���Nf�L'�r�v���X�����c�:�����l$�CC�Æ�2��*_�����󗚋�l���52��՝�I�?C�T$(K/�=�נ����>_$�IiW�p;5x�p���uz)~Fn�,�Ufd1�3�;���^�P�vX���&O!v���0^[����2�If�o��7}J��{s
La�Bn��Е)�se�N}�/K�j��(�����ꎽW�d��<mȊ�첮��^��`X�Ȉ��J�gd�z�=+��_3g�`�mظz1bH
_;R�p��k��z�%�<Ͻ��r�z���R��s1͏d��ρ�:\W�r2���fr<Q����O��k"U����-�.�}r�}S�P�Ӎ� Ww�.��=\�]�Ov������g���@�i�XR����FW`����v�GM!�o�/��t݆u� >}X:#6;>�HuyN�6!���eq(��?X�@��ںZi����]�vB�����Τ�{�e��꒶+�8�ap���^O��Wɏ�
���j�8�X@p�Щ][�v�u��mk7a�[��%c�7s���2��^/�<���w@�3�y}�B�����{%bʏ�Q��Q�{Y����Q+��8���Y3�\i��<t��E��|�v�����&�#%�d/�0�FUg�K-��u�nwj����ú�yBs�}eK����z^o�����������[X�e+�����*$1�$�k�L3�������Bxgjkso�"���$�QW5`�-)�7�A{�G'>* y���~�~�����ܒ�=l�2��je���HEDl���Y:�s�.9�~�>2`����s�y���v��f��!(�f���F7F�CO��L��cd�Pr�@BxT��� ����Q���R�ņ�Fi�KS苌"��d��G�ۅ�I���?��0u�JS�̐ʅ�����5��}�op��@����()n����{��`Ԣa"���tnu'{~�
��;�����"�SN6(TSi�����`p[�20�����Zy9��zX���4@�wRM �xr�'Ce
oy)j�mC�Dl���FS��>x��8m>Q'k�qzZB���q3�;��D�ӱ�}������M�Dە��q�������C�L�~5e������
�9�[E�����a7��M���?[������Ko��Ό�(��} S�|wB����ܴ��m}F�|�Y�2cr���.(�
�d�0�,Z�ԧ˷u�	i�-��۵�;7���dڈ�d.nŉ��q�5�nx(3=rg\�ީD6���ᖇ��g
Ra]����G��_e��H�=θ�a�n�g��c�b��:��pUr吪T��W�^�N����r����	��7H������Α��A�]Ο��e[�XY%��魥��$��.�~��j�ݰ@9�k�|d�2[!:�U�yb��D��^ߴm�k������C2���2Dc�	x�0�������AL��,�}�Z|2�h�=h�w�XS���5D�ٔ���.��!���z��bD��DGuk"�F��>*�>kC�r!h9.�q�7Xd�)Jzf�'�q�;��jA���PT� H+K��/�=�l}ݾ]�鉡�3�'�Q�un�a:aH�����r���E����6æT8�?�`����X���9nvΌ�����vM�;LR���mTH����pJEf�����AnO:W�+�Kخj� '���|��;?�^��\��2��/�B&����&`}�5dم��#����Gֲ�Ø���g6�E�~��w�h���Z�.˰�K�����,�N��u��Bʎ���-�j�Vm�p�M7+Q��r�\��s�9��\�2C�*P��ִ��\��QG��OSQG��v���ǘ�F`���T�=4Wi=O`ׇ��&�����0u'��xq�؍��r�|h>b'LGڨZ�B�? ����8��k�$��(Ji�V���Lo~0��b%$� u)
��/��#�P]F�N�0�͵���0R�HoJ�d$�t�Z���2�擀ma=;�3��2%����yvVCD"���N��߀4ᮼ-(��iˉ�R���\9�DW�/D���m>l�h�v�ى
��{�t2��3�%&�c�?>m�/rMC�P��H$^"�X�hpxѢ]�:2��#���c��}�U�L�*
v��1�R(�H���/������@�I�wKV�0�zʤ)�Pc�G�8|O��Q��l[��bD^����[�E�a$�z���^7t3zŀ�)��(\VДb��@���v�P�*��8𭺣�I�BD�I�޿�B���n�֥�Hto(�[Hi�E>���jL1��	F8���4aH7����f6�Cd�����.���'*hN�ST�5�T���+��Ky���59��4V�+�o���P����C���w[��e�ڕEE��$f��\v$<��/�����@�7�;�F���C0�b�W��Sp/di�p��Gb��^��$g�WiE3o��s��){r�@�q$q�N�f�����X6<�9X��GRL�Z�I�vo����Q��H���z0.�?��i�(��Z���1kH�î	I��&��.Adcl@��[4��I�Tr���q�cV���&�(���>�.:ma�#k���ҝn�?�e��R����͙`��1х)�4 �T�F���7Zw��nw��F�8xq���G<��<B��Y�隫��O�"���#m�E�o�K���Ta���üO�)��L������GH=�C>�9�\[�^v������|���12������4�Y5�@]���M��+hK�x�~�H��;�?��5E]�<��;���#��k����͂�.שe�I�1fvA�Dk9g;?��h�m�>�rv�T'f2B�+U[��@�:T�WLW��z^�=�,�K���x�۲�8Fw�7-=*�\�:p.�(��������W���>0��HW�(�v�0@�Tql���`�:W��6�����2���.���
�T���E1Q06�>pJTH�d�
f��'Z���I�,���w��K�?�ۋm¢Xi|��r��G�8L���g..Y��EP,��2+�:.&�T�`��������x8t@���u�)Xf'@�.7@��'Vi@^�Da�Y���Ҷ���*(1;�(�_�=����SZ6hc
׈ k�G9[��W�Z]�n����A�c80������v���G����{���4�Ќ� d����jۢ��rk܄d���=!`�0��ɵ6�X.&�U0]q����02�/GP�C�g��ʥ��5�;8��\�8�Y���1C�i�]1�N
�c���u���ӱ����o�a{g��5$��^���J���hgU���0`���29������gM�3�D�:���F{x��1��� ��0�e���!״����Cr��Q&� �,����=�ǧˠ�a��q�仵2&_��t���-�Z�y�y˘���f&l{��3	d�*��&32�-��R�(R������U�n-Lo�֦�C˨@c氪�;�W��7Ok]�_tS!q%'���(��[#U ����im��c|F�	p|��q����2��P��>{=�u�,4������J[>�+]:j���P/�4�$���8�ҵX�<�+����{�`�6�P���p.����.�m��V�#���:U��Q�^}��4�p��>3W���.B��]6���^TS�A��ꘛ���)&]1���Z(��Ռ����
S(,CE��E���-�z�,'��Ɩ$��b�ɵ�����~�@��r��\�WN��|�*ܩ)�;J�H��,��?�]d��t|����D��3h:<Đ�QL��Ρ�Y�K����2��|�m��#m�@S�!O7�4�K��<�\g���<~�W8�ػ��t�Ŧѫ�����+k�h��mŦ�O��ȧ������ �����eτ��Oz�S����a��&ag�Z^��U��Q��<C���R��sj�q�,�a�gGNg($��;8�mz��ޣ̚�
q�$��t�^c/���	��L��Ȭ��F���ҽ�W�ɕ��u���[�ý�0m,`�uh~Yv��©��C����&�Dݹ�����h�g`~]"�ٹ~C}[�:kŗ���kE����M��222yRP�1�����57~��gz��8x�]0�l�U���b!����-�/W�$��e���S��B��$�|���u&�tUMc>��]p��L���z
b+��N�ĵ�4w>Q�*�������}����je�L�}�f��!�|�7�O��I�e�%9U����!u���D��vE^�d7���*E;���CQ8�u��+Kt�M'�����M���2 >.�e���=?�����韛l��Mi"��t���}K�9-b�F~^�7p��6e���ڿ��^B9L�m/�����O^of��?o�.�\,���QT�����*e*KM�ˎ���ˈr�Ja�y2���ph�=���|ъ�wJZ�������L:�nR�����z`oݍw����/9�v�`�Tg��3\KĽ��Z|����I»��c�w�ҷ���7�a�p�M.��VR�Xл���sj�K0�b��貉��N�߹���d�^v��ɨ6؟�
T+��ʏ;O�\���GM��.�ڍi<$)��P_`��щ�s#��`� T�JW�\���;#�C�Kq�j"`����|����c��ʬf>�'��ŵ6l��*����W<5s�<�����w�v��p��85���D�����@i%�x��R��Fh:u���f�WFǲxȟ��b��ȉ�x]v���'3�U9�=��l� �+�E����po����H��M����8�O����I�� �|��������T,��.�*qqz&��d�6�����rj�D�5�
���m�`��g�#��l��+؏^�u�t��s��ʤ	���*o�X�Y�{�Kx�oxlWb0w��y&O�-]s�DuYިh�Qvؖg���ѹ(W����pRSs�j��m�!<^N0Ay���.mfPY1~�"Ұ�۟O^ˢ�?�ϧ_M(],��q��8����iSwl����A�H�E����q��y�ɑpz.+~���a��c�UM<&�|���?"x�.N���K��5ɳ���B[�8*��k�
�Q�}j��B$HO��6�9�6cӬǯް��U_ﾜ$q��5^NY�&��Y���DdI�1��t���vo�12v[��h(<Xx��Y����-�V�PBn���b�x�
!�
a	̆`�}@t��f*�7�s>V՘3�O�e�<':Xej��ύZ��#[����(l_�b��X��l��ڊnZ-0�5?�INh%�_�	����z((������ �;�d�7���|)'q���H��U}��|4�C�����0�3��=�ɑ�Q�q�M�C�K'Q±|�˜h���&��L�R�ˬ`���x�bVĀ5D��1�u��|�D�H7�E'��|4�����0U�=S�I���@~��-��������~�$��r�S⴪--�+��T(��e��Ѧ	���ez˼��m���p.�7�����ͺA�؞w�g&̏��*�w٫�QOTo�������Ә}�3QɗN�4����[�߳h��>��� ����;����[(MU	V?�d��"�Z۶�j7�P����]����	1��;��+����m;���aNQ��=`���mOH��$�WU���ԑ+}~�싍� �x�ܭ<F�1����w�O3H��uOm��J�wb�8,D`�^兎 �IK�2��^�	w(G�+E�W��p&�F]���I<w��N�;a`��X ��7��+�(j��������9�p27��j�f^]�*ЖU��!�7��f-ײhz�/�3��6H^��a�5nǨ�}ҭGc$��K�׬�A�� rh�.�&���z`-��tێ��Aa+�A���z)rD�%��h#�ĖK!��>���zG��8T��;��Scj�	�6,�]�n��R�F��F$7g��$-o�/��t�V�/���1n��w ��Kp���������D&�45�x�H{p���S���ݴ�r0�@�~^L��(S� �M���z�f�������@��n ��c4��N+ Y�y�*�	C�8�c/J�#�� �(N��
a7o}�l�����Ei���$1�!Q�m�v(N����֏��5�>�/0�e9Fъ��+����m��}R�0�Q�^U���Y�ߊj���g�a�A��T��������A�&�d�l���>�o��P��y�b�G⥃3���r0����:�mm�Z�ׇ�9�а�+b�	�t�s���[�l�D�6�Im�Bի}�aPX6�g�v��*2�'�X�'�	�܁˥S�>����U�%����1o��M�=A�K��������X��&?��=_���=��t��B7x/i�Ȝ���Q��K��8C��5��C+����~Gvan�a���f�f�������6?j�f^�� ��h����o!�֕�n�T9��V�w�RN������T瀗]�~�[A`��P�}�����w ���L���&TQ��^��U���i\�}��A�V��*U��<x������V�d�������yn+W���L��}�X� �� �Y1K�&�-��TS�hp�|մ|m�;��\�ok*}�}c��b��t�)�����M�ڳ���R�5�i��)�Q�����Ѽ#�A�o��B�6������"����n����^�;R*��,�j����h�ΡID�kZKZP����n�|�2�<��,Տ������:h�互��FL��T�jI�,����Z#����X�l�n�7�l4E��3��):�U��eG| �;���/թ^�¦�{�*+ls�%:ם2�
�V07�1�J><��x��|� S-Laӥ�p
�d�fgFj	�,J�P��Vt��1�j��D]���]tgj���wt摒�Ǧ�9� wMK����U�:-����ic,M�7c�7:f��=�A�5��\O�zt��+�
"�ʾ+H��u� �1�5R<eC�*�5�t��	:��~s�ez�򖃤�^���1E/Z�����v]�j�����Xa�![W�Hy�>5��L.�#�X��[�n8�[���y	��/`�+�Q�4!�`��(]��+�jU�e�Idƌ�
�zu,�Ǥߥ���%�P����n�;{��r��V�#��t��;��/
4d��_C�U��'{�gZ���o$"��!���'����{j�Xuđ �:Bu0�a��x���h2�˸��^�KăF��?�f/g�/Vx]�S_�Ls β&���e�I���1���bH�]3��x�>�9�m��.����*���A_�W=����Z�W��U����<���J�XN�A���s0���s��$�����|D�4�	��Tڽ�uzn���y�ۻ�_��l\��k�g8�ۑ4�	�!]'g��4�#��i �|��������*��r���F@'t2�'C���#�Q�����C3w>l�XDՕo�x��Rs���G�qQ��O�6vu�h2�LPb�Kw�7�}�M�yV�R70�bb��d����f#@��ĻEA����R��"^���2��)�L�y��/��|~c��H�~W�F��U?��*Xڡ����A�~������2����Aؓ쏍���:���)gn�����-�1՘Q�H5x���K)cƸC���'>h�>��L����y�آ��3��b�����d�©��R��p�:��!
]xA�t��˼�q�-�(�Rƪ()��.Υ	"�(|>�<�c��Y��It����Y�U��F�H�핇����Oqa����.��!�TG�/a^�l��K͠	�	��L�L�o+�o��w���=e���:p@އf-͕�$b�{�z�j��(�~y���3�K��OÕ��$b_6^�L�,�@RLB5t�Gg�'Hɫ2g'oP��m�b���C�����C��s��:_�q��+�C?��2f�b�}R�z���� k̢pR�]���ECb�'(�{�ޭ�~��j�v��+�����|x!��ÞA���|��7	p���� j���ǩ�J��:U��3�`����Y�Esf����ןۖ�J�����9�a;��A�- t�և��k�*�e%0Ԣ]����2sު��ע�8O��vY�y^܉�����$(©��X�Y�j|�$~y)���`�t�.���aj!�@Yռ��� C�9���;�1��oE,u_U�S���6r@gѤ�ɬX�5�C��Nl��z��gI[)�NhE,fz�R��~����UGty��Z^�G��=&� OY?��S7
�̫�p���&��>M&�gE���,a�$t�B桼Q|�]+��.�8�R� �����اm����\��9��p�
?�F^f
����&�z�~��� ؈}�!5��������)��F~�:�f�� ����2]D�g�dP՚�]2�ԃ-����M����4�HY�t�0 �fN�^rT��m�U��9zBX�.Io�o��+���{��0��A#8�����~M������l�O䯿��V<������}}���5R��Fs�Aa�9�����[�D�ЦJ���S���=�;AO�
���[���d�°�vd�;����e�2�T�8_�	D`W�e�_5��}h/
%�T!ՙk[-RR�txJ_`��N)�N	w��U4߬8���Ʀ�I��&y�Ut�AMD6pl?��My'���������
���Q�֍�w��3M� /ڱ��|�[��(~S#�_�v���9��$�X*A���{�������K:�%��Ui��;�zA�̔��M^�%���d'u
���i�n�^�=rr�}���j,}��O���>�X"aФOL ʞ���`�uDY��j��d�3��?ѡ�B����d�R�&�����>�m�&�ו4���i�6��i�R,_�u�_'���Hnǉd<�o���ĜH�A��fl������z,H1)i(<J
�,}��Y��4Gت�D~�u�FO�xs��h�u��򂥳D��~7?�?�o��C��$g�r�[d��z�J�x���fA45o��~H�>���>��w9
-0�hj'p����E��S����O+P�>�^����{�����rp�USn.����������X��赵f�B��NE�@k+��LNt�̺W;Jc�}.����x�_���ԝ%Y|r�ne��S '���g.�G�\��_[xȰ������DB�&�U�P���:v^Xp���`Q54
(��ǭ��R��9(ǈ�s���ϋ��7Y�7 8vӹ<�NnY���}^y40
jì%���}�>��I�'�B�x�
g���������UR�4�q�T���>�NV�ٶ��^f�E/�܌P�\���� ������
!2���#�u�5�������7�P�?KV$���E�KDSƧ#�����⠨�!Z�xKI��c��1Qd��*Dk�,O��]�V��vn��	�������^�6�Ty��:��0��K����|dDq�{k4~��7�S�MS�W�)��+}�B/J�~���ܴ^(}�����K]���'J��:��f}�@�?ߐN(�[�K��D�-�i��v�80Qtҕ�(L�63�a4om�2N�u��bp*6�P��[i��e;^R���`���j DCpM��j��9�0t�M��R2.6J���j�B�j�u#�"*%��΍�-a*��f�P��H�;��f�6��d����B�$>g���˻��K]x�Q�!W��b��`m悿��
Վ�o�5�`c���#�ã2�������L�&��~d�`%l�D1צ^��PY�d�N���~[�?e��	X#��cqh-�g,r�_����tb�I}EֆPk�[.�`�-����2\\J|ࡒ����tM'�Ϝg�ww��K��hl3
�v?���R�y�7�0GI�>	�0f�� K�tї��}]��},�u�9Llq{�&��GPi�V�����g�g�Qp��=f�����U}N��7�����̆Ԝ׍\m����E�O���(�*����ĸ�Ʃ��C�Α!���\p�w����d�֭
�T��W� ��`d��t#W�OC<��F��@N\pj�$y?lݡE����њ�s���2��mTm��vc�_;=��fT=k:q��P�����G_G:JP:!N�Y��g��m3��UKj���U)�'6�4�d��[5%�`�	�j�U���{29�� ��W��g#�h��&OD�O�Îh6f�����xs��5����m��'�\����,����Q�������S�s|s����� E�	Q��=s}�"��r|��.�[ba��%�	�=�-���6�X��tp'4*ط���з��MT\�Q�1>�\�O�\�L��$��+bv���Fr{E��Q��\��؁�e��W�C��C	j�vE�a�2/�c9I{G�`���X��K��u��T��_��o��cd���>Z�S�\�ݮ�Ѻe��9�Wq��xH9A���_��]V�'r|�4��@�a���	�?����,�(��T�UQ_�'Lu޳��*^���,Г��!Nc�h/ݏ��*�+�d�lƴ@E���n�@�ߚ����3��S	���d�$�ؐ��8�7���gm�*��œ�-�>�H&�}ۯ���NVK�4��~�!S��ߩPIy��C�}(�f�$��z��2=�M��sc0Hy�d����� �L�����ߌC4���#�9 ]�ӡ�Kx�j��D�G��[7���e��͘�� _�
7�F�mb<ۑĿS�o��lJ^@w0�y�熮砾A��Έ��qP�s���"{��=x~쫋���dR� ���}&@�G�T�ݎ������-����V�|���̇đц�lH���[�y����|;�4'�)^v-�������� E���/�[Ӊ��ƺy�g鮊�l��l�������J�	��$%F���9��C˾F,5K�ۈ�0"����k�HzG�o<��@]=��|z%���l��z�O��c!��~3l������ ��,Ĕ�A�w��R�܈�:��LP�?��u�%�jWlEr��"R�����@7E��O�vp�֐ؕ�o����N-Gs ��l�k�-v_���dU WJ�g�{���e�n�G���΍��|0S*���,\�S\�O\.ɸ�]��)H��>�6�o�!�}v�sVdY8��L\	 ;"���%��2+��� ��XCQ{U� ����v�XV�/�Y��-5�gL�
�]k��w7���}��;��D��� h�$��.��6�c�ਗ਼e��
�UP|��R_�B�����k���W���Z��'!�3�!S���r��Ϲc�BH�j�R���Ȗ�c�N�렄� �h��T�����5����P;ݙ�Fn�%d��7F��걜����h1NY��!��w�e�~
Q71�*;OW������S�x?��o�^���]���\{wo�\+-�d;�g��D�3�l@� yu�ŠE��o.z��Lh׶鬙Y@���=l@Q���O]2��T�;~H����.�yU�i�����-��ID�Ћ*'#�M��U92��c.$�������X��J�·)P�lQ>��b!/�Ĉ�.�<�����qV��` X�At�`�X\��"�����\��(�	� ��ƚ��9���lN�~���f�F�?���~G<��k�}�5�0��J��?��0R�:����,�c�[Y�M�mB�9���|E�I*��º�o�֙ a~�
�)��B�e�����ՍM\v�~��30	TD�M҄���)�t. �D�Q㮹������Q����*d�k�>�B�F8��oZ\a���cl��3���c�E����卒�֩�{�D=Q�n /)�>� Mw�O�A�):��{'(!<�N��3��/����ər�	I�&�&�#8����P��f�&�MH!E�@�9Id]:�������8k}���ǎM{j�����BS�fd�*~�z4���I">�� �G�3�:[����lw���K.�R_�ޅ�{)x}�T�0��i]�x D][�u],��NDό-�b��E��$����� �pQ�MY��]_��`]o!HD�w��\��>(Y7��nS�-Ie��!Xel�!0���+�@����fP�]��9���&+�XB�N�9�
�C��� ���$���D�hO�P��r�u�9Ǌ�.���2�	n=��e{���6������*n����hEU��:���V���}@�I�q���h�/.zމݦ\�C��z$:6A�2ҩmKC �RB7B���$�4;ޚ��	�a�>	ׇ���L�!��p8K4�}�õ�دw���,Ы�����2��_� �hܵ5a"$��E%��v�+e��a�r�&!�Q�>���:E��jN��~�����9l�HEֵ�9������>5�W�D>��h�����������G2�>� |�a�1	P��]���#���=����
�t#���s��F�^�+q/Q%yS���IH�b��������T9�X�|Aó|��t��ZOި �S�O$U%Բ|�	E��%�Ϭ� 0/�_1�������jn4�P�d�G�@��9���t'�Bb
�O�q�&3���1��W��M��K�\������]���-�CQ��B��Dϗݩ|R�
�>(�#6�1$Bo{�>A��6=�pK������V���{���0?LM�!&�G�)�:�$�4
`X�<J���Y�"oﳤ������@�+�=Ek�&����f�h3Wm֩�@a������D��s�
b_���z�����n�őFg��J��p6���R��Wۡ�X��Z_gl�wQ����ϓ�k��8m+!�)F����^s/9�jda�sym#��i,�9�DWc�.0p��t���o�����1��Od�~ ��鸙.�zxm�p�Զ��e)mG��#�����9n��I7	�J�Gc���dg�H�6������)�	F�m�������m|&�M7��S`�A�˨˘��c�����>Ӆ<�4٧ц�!b�f	��׶B���ʔ���	��7��tM*vs۬�2!�O��c�0�ud�+Ck(Z��#+t���_�����u-�1o�:VCI�b����)rɎ�ajG��*����pځ�>֤+��t*<�&l��E�.�_5����+�	1�'��8����[����V�tM���́�v8@��i�펞���@�R?�U(P�9O��)$<�,�M��N������g�.��%K�$)u���T�ׁN����ŨZ��RY�w�k�͋�>s�<������f�,���M-Y��ӑ���~ۙ\��>�^}�v�n��Zl�)Pp��\Ev���g,�u��K�gS5�R"�>dz�@�U����Q�Y��L�@�ߗ �dr�pL-�§��X���n�ۊ���`�bY��޾�D�����X����D��t�b�-B�1�˄�f�I��.J���o�T����Ww���m$�-�����!}��p������5�pKzojsS�EP���(�j"�iv��/�F+ð����p~�$ �h抴�]��I��C8��A�D&d�DO$��9bG�ɐ�}�x����:]h�I,�����G�?�m}T�N�s
fgr�;�T�e�o'R��)��>\&�����˯y���F��P$d6�4�K�|�BЈ9.wf�����
�tw�!�ĂhJ�:t��'����_�4KNU3H@g�Q����\����0�ss�Ӡ)��f,�C��w�Q�`��&�N%�Z���-���U|1�-(Óݻ���B��\U$D��{)�5���C�y{�cQ^�r���ڬ�h��D��P��	�^|qh�����L��V>fQˠk�� �D>��w
M��UL��o�}��:X�N�W�/��JҮ�=�a��y�Nhϑ�=���9T�[�p�*4����[MZ�bw�	��M�4W�u��í�?Pt(B)t�Uk%��\��P�D�P�r"+��9��ɗd��_DjӱJ�]o�h�	/*�6룏LS5W�
GN �R���A���f#���}(Zr݋�;F~#(
�������%:��1��e����{�[��rj��"R\%w�R��sJv�P�i��\4��
KUG��:��&�[k#r~f�y�B�L,s�]�ԧ �O7���-~�CL`�6e(P2�p�t>��� D�#�hZ����K�v�Ͼ5<��:B3+���b��r*���IGle��V�ڬȨ��/�	���������tX�jJ���l��g	�d��L��!�(�a�U'�x'V.�p?� ��$�`3����-�W?"��U��H��+ɚrbI��Ӆ��1��l �Z��kvm�1�%6d��1��_AV6�\$Ofe�Xm��:�gSf��X���{|�n��1mh�~�w����Qt�RE_�X�K>�s)����F�jW�[(������
2�%+U��yB0�+�{�$4^��s�w�`3K1w���ą�}
�q�"���5���jfQ�����j��C��]=���*	JY1�'3� �G�<C˿�?
0d�t#߈�lq�l�/�����#����ٺ�w3����R��B��e��}�q�f�6���g%&s��B\�>P֦���h��V����?�A�(7�F��v���\��_��H�ң9@^�?f�	�t��Y�Q��@��U�In���! /��bX��	݋
lhT�]|�6�*y+U���
����<l_8_��B �{�yO㢏~>�6>A1�9)�@:�&nR�c���Q#_��D�p����C���� �rj8pm��A3�m#A�0g�����z�Z:@�I�J��-�}� �՟QF��o-�Gzѩ;?���g�Y�ף�Rt������RZ�a�𡣘U��b6������!$����ͣ�_�#� J�XZT=t�y�$��.B������F��!��6=�L��kp(0��Ō�$4�fa����h�,5�7�▀f���z���Ҽ#�� tA�Z�oWH��hj#u6��(V�D�9	��,X]_m�P7� Lf��if	�J� ��ğ+��y��S�x�����Z��s!VamV��z"��>J̛BC��ى%ղ�m���'�:�3gk4��N<���
�M�v@�����#�!Sn�aM}U � �P�������񕻿��Z[%����.u-�5p�a,�T;%���h�}
�,m�[ Y`�%���t>lN?-.��RJ�a��x!�w�?���u����1>�]��l܄�|����6�6������ۗ��-I�p�U��Dvh*G�~�v��B��Z��SRhRY�:2H�ա�Y�9Lm�z��[J�Fʑ�Y�!܋9ޞ�9)|�:��uW
>M������7��{�����5��������N���>�	K��֊���Uz��1��l�:�,�� �	 &RO�>�x~�]]�K,}�5Q���CC�g��"�=������ǳHW���E�=$t�J}�&��z����%�g��F��.�`��89��K��C�)��d-M�N\���*��&����9�̚���֥T�8Ǜ$��\ea�y���>���5\#�.����4:�*!�t=�م���C����g�c�o@{�u:�4�)IE�s/Ll�;,�-.��[��wm���[�#���o��6a,<�<��vǱ�9�#��]`	W��/�v�	��e��C��p��z���&fjz�u��J��z��]�ˑ9C�ۛ䣾���%:b��!;�Cc�r���M� 6!�(8�mBN�!�.&�+����6�\Z��d��J]qP�M�(4�;��3�ܹ��9�WFNG-t6�G�Ӑ��R�5G�Xr0�z���/��f�����ik��J�@�==]x"!pZ$��&O�?�{wp��|+_��)����rY�ѮU3˘�'�M����
��rjі:�ͮ��U	_���:����6\�/���ۊ�g&�c�V�W�O�n�I8d|�pP)L���?J�E%.^(�A /^��JS�d�hg��Oa���`�0�۽�gLpo3�����#��}N8�W� � PV�L8��E(l@�-#q�ˀ0q����w�T��v6C�bJF��:I��P��U�v��	G���JW��!̔���	�Z�x&p���zԜ���K����$��Z�J�N7Sw��0`�1����AC�0ϴgVk%�th1C��������<�G�N�� ��d@E�N�~(���<�dİ[}�~��ͦVp�5j@�����%7&�C�#KC��4�������1 -?i� :�����q���{�M.�uU1�.��٣�%	Q�	�������cpW!0S���U�����t�M]�9�P��?#��.�����a��e��Ҵ���	=�&+f���@,�(��QŽ�f�B��hT�Ř���U�*�R{գ�^��t}  ".U5��m��OP��>�8�t�s�}�IP3�o������{�% ���/���P�bv���	i�3f�Rw�d�eR L�E�#�V
d�u��!�D2�,%�и`�ю�K�*�%x0"k�0lC���hJ����Ht�4�7�%i��T�Rc܍K�Ѥ� у�':�J��d��*J��x4Π��M�F%�A�VG�i��p
���(رY�M�W:��'[9ʭWw̭�

�� BC )j�K;��鯼�5ɨ�d��2�ka_'��XPi�EB��~���J�>om!�h���vg��4W������D��Xa��S��G�J��o4� h7�H ��8�C�d�x�Au!��OS�4�m�ty�w���I�����U*/Q����djܡ�}��ڜ�r�]�(�?I0�]���՘�1�l�aԉ'}��3{�Co�_m�7g�	��5j�
ͳ)T��1����hS�&�`>������=�z�St�9���x�&r�B�xM��͓ ���BU�mO��KzQSz����1ܶ
�����������rF�����wVH���Y���]�I����dn�� 5��~fAl]x3�,b�č�@9AXȞ��~�ḓ2e�>E�=�`[�Bqp����7�����}���β��]��\x�r�#���敱%ο��C]�#P�T��k�a����r�)̄/�`YiC�3O)���<"9=�އ�Y<���ɷhT��՛�n�:�4�.�]m�͐�{�Qת��*�Ykkoim��󧉐�朅�&�+�a?��o
�4�	���i���^P��B�NA�2Q���(�ǀ|��8δj���81�!6J�ֵ�&L}?�UQs_{K�o���6��B���tj��6�;_��%N:\�&��~#�� ;#�>�Kj��6!��t�=��Q[��GO����e6n~-�=�y�΄!	�C2��������f*)^����$����-�6+�X
�c*�D��46�恋?�s.I�#N,g��Jwvu�'�<�	f.�ӬI��ի0Lʚ}��.���J��«��5#C�ѿ�'�1N$��)�а9�q����b�S!��xj�Q��y��n�W$����
U�TFk�;R	�CT*�ɉT���/v�3��!�e�c�����jh���E�
�rs�%&M������fc�<�S�6w���D��R����<w��lVQ��dGBw��x��Χ*�2���t/���򇃟��?V�|������h�,	&��;A�duF��z�xЖA��ޔHb#����Z���4U��}
j���zA�՘��ˍ��t�4�������Xt��ڟ��KΪ^��.\�,�N}�
֨w�4��ޖ>�ɂ\�(8|����GK�%g��!�<~��ep�����x�\$��Ƕ���,t\��x:��P?�zZbJ%C���8bԯ���8�����{�S1�4� �_'h#7�ѓ�5%+r�*1)�o�p�T���WB������jQ�M+�#`�3�aZ.�E����.����q�Y�OГ'��.+�U�z���N=$��M����$�s�Ȗ�Q��w0Q��b��^&�-�Ξ,aA��6�Gb��e��1�w���Ȱ�7t8E������m��pvs9�J�g�]��zz	B���3q�@��D8z��N�Z'�0��[>Š>&$@��_C�|��]��E�%^��g�3 �y�ȱ��;Q����jD�����wtJj[��$̯�{U�ʵ�����]D�-0��	���4B�B찺ݴA%ҋLE�EL@BJ�-R���n v� 0��.�I�e��[{�L�x��a�� 4��WW�V@ȰuN��矃��ƙψ>j1��G��j�����]k��Ҫ;|�%�6B ���$Ƈ�GD?:����ڕb痐�/_��:���0��>樵k1^kǼ���r*}�Zq�2X.�,�+\es�Bz�?��.^]���D��KCdH���и��3RY��D�}#r����&�/uYx���e4�t��F����S5��v����}ҹ��,[�O��y��7.w-��,��\��6��H<�g*1b/t�]a;�X��cn�70UT��c�����c�A`�2�u˽��W���r�Rx�݄���0�T�KM�,gG(�!�������B�|b��xcy-��%N�
:�2��,���ނ�4�B���M��`����s��]��6��0+iy�@���aHb��8�l@�L%�w��2fW��S|�҃a 'i���7 ��T@��Q2���.2�"¨�r������qy��*�B��T�)Web&9؜�ݪt��쨤|Y#�g�TN����Ѵ�D7�Y�m���~Z_�0D?�O�ׂan�;ۯA�����:��>�A�Ot\T��U�=�?U(C%)��4�P6%���P)�;f��+U�����L18H�e��\�
�d�Lj`�a#h5��sC^�Fg>X�����AE"A�r���G�����Ǚģ0��Ȭi�q�Sצ�В T�n�(ܭ��ZN�v�8"�a�1{��n�@�#G@���`���j���1���R$���ݪ�gS�rpbg��H9iڦՐ�jYc�n
=�tsC����.�>�co"\��Z�(lV�L���3e�R��|��s�i5�&xZ�I��y��K�� ��gSHn�'ݔe�eM����Y� �`�&�R�Y1��rV�7�����nF˫��·�r6�2Qџ/��WYYR{؀S�GI���\M1�n5Pe͚~�l<?Ѝ�:�͟�1G^\��EY<._sT�PM3�˨\>"�.�*���9�j}?^0����{_Y��rɒ}jL�����[�/� MI���������:�hig}K2N/l��ȋ�������)�EiC���8/R�<�yj��F��l��k�vg���=���j	�5�ѿ3ssD�E��-~�
����,ŀ�Ye�FH+�K����Df��ިd��Q�	�\�F	E� =>Z5+�/��KڼM�v<�G�c ��R�|P�e�ca�H��3X����)�Қ/^}��C}�3�n��Sz���`nE�B�A�m�Wj͓�YHL��z�Fq�`��:�l�����6$�).�u��\��Ü�=�2nj�VD��]Q��T�����w>{�_	p�cQ'v��.,i�@��,;x����vL�E1a���]���l�15��x$�;g�Ԏ=�ܕp�Ϳ����7^53�_н�����sS�� �cz-"h���nU��
��m��4:f*t?�%#uH焱�:r�e�L�\nU���v�`QQ���F�ţ[l�=���y����mi��F�
s�D�V|f�Rj����k֜D(��	����&���Ql��K*L�uGiQ��I��C�m�I?n��3�p�>�����������TZ���Pv
�u>=���0������w�"?;�i��U����03��Y�Ԍ]���^�������`d�CT��u��4�E'5�[��b�`��R~b_��Wp_��`$��Zǵ�f����$����V|�,�Ș0���DT���":<Y��썮ΐI��������&��^6y����)m
���օ\�r5�q7�C�̩�n��#�Un��vf�ؖg�| �3��bp��pm�sZEч��+u�/�@f9���M� {(�_��Ι*ۤ�����%��:�jI~�'���N�����N`Ԗ�)&�sp5%!�*Y��9pn@^Dכ�ҏ��ͼ)辟�G����2��Sdcq
��pu3gJ{�%k��	X�����/G�$A�7����Un�S�����d�S$ƭy��Ө��7:^���
�0R%�G�07V��rd���cD�g��#~��d�lqQ�Y���+]��YF!3�d?_�~�&�~��ϙ+ �>�n�䅧_��P�W���
e�6�E�5�e�ޚ�6N���."��%MRG�r4{�V�φ��,9վ�
���AϸY�bǋ�%���@��s��B'�}�T'e�*D�I�`��٘���O]ÜW���М"B1�qd�BQ&�#�W��g'Ty,�5a��!Fgn�NQ�,-�`f��o�?BY+\�#��V� \�~k�O��$gM���4�_� ��qfsh�rY���(��H4CBE\�35���k�Y�ǋ"�����v���a��,!�/��ے��(����N��E2�«Ղ&���}��!�s�+O����)vH�!H��K,��L�&q��N��E	�5�b���f�{���4�r�N���M���ؼ����d�w����9	�����E@��S	��fs%x�P2���Z>�&���x6�}[:)��j�lJ�Ғ{�M�"�=����U�V�Gִ[e�t}�)��ׇku��ق���g�O'0��4e�HK�{�GKѢ>|������ۥ�oc`N��� ����Me�-�OE�����n�a�����~��3,�7�Jٚ����p]՗l�-�D�F�����{�wW�C�Pֵ-l�{٠�4˾q�Y���t!����Rn~ϝ���N��l#��eG�S��"�:�T��N��V׵�����CWO��m�>Bi����3}�b�Co��6����)&���jw=��Ġ\1��67�5HG-�n�9���j�8��ї����ip۝ZkP�.���$�A각p�p�G�fE�:��#�G��)Ȝ���f4��:�2Po��CW���`�	&?f�$d	'h��b�Ǳ;��f�o��j�"��Km�K_�Rl���$��b�\�Z��;����iN7),c�~w肓�\�1�C3[Y�R��L#>\)�>�.nԵ� Y��]�eT�>�D���� XLu9�M5x��p!�RW�⚛�^�^zךbq��K	Z��^����|���;���G4�Md�f����k�Z�[����u�@�M�N屶t5\�J�	WS�qW3\d�.�O,YU�����@5��(�� �t!�Π����}��I�T�` �m��u`p���#���Ø����V�%	�(����1�<�����?S#�9C|�L�i]��c�_�SaB�2y�#�DQOD��+�ogܬ��ػ�"�I�Fs7�{c����4����4$Q԰�k/�Du�����d�n��K����I������EĞ���z�%�|��*h���>4�ی)�UҜj�N(-�eqG��B)�@��?�����ZA#� s�)���� �PMQ[�������uד� ���9����Sr�w��~K��Z���e�Y�2�W���Z���{�1����6��D'^�'oif�������>�I�dt�20!�V�����O����LZoO<Eq�����f9����ѵO����4^�!$
��4�L�e��_(����Rǎy�L~�y��:�����Z�<�s�}��/i=b6w�b�o��:]Z��6�Y1��X7d�KH��6ސ�£�����,o��.�$<� k�f�LY>��k���;�"�ɞ�F�r©�@:����k�v*}����"�F�ʡ�N]��p�����$Z�e����$�m�i������>��Z� �=�l�r��QO6�]����w�eZ��we^ѹ�ޠM��!j���B�R�v�a<J�a���)nI���8��d���ù���ͥ�AG�w�X����O��)�2K릦YO'�<�9&%���S5�"���.��l?��lm�wb��Ubޗ�����Ѣ���;�8n/�4Қ�-�`䃪�t�a�E��&�!��>e�6e�}_�彗%�Yx���9z��R&|��v�(��s�A��:��xR�KZ��%�h�0������<�J�%ZC�Udi�]�dh`H�0���H�8���c��;�M�pt�������ć�{V���g��t�;��U��f�@���
0HVo��%Nu����h���p�`Oy8�����f\��J��=���ԜX$[ �g�/�sC���r�ADg�i#��̶�%S�K�TM-�ڟ����	�r��kZ����p������H>��rC�b�g�
�F�����|]���{;� �������0��NK�*����ɧ��T�C9�����za��h5�E|,1�b�K*�]iʐ�m��8�|�V�$� �9V�������|:8�ȥ3F)�D���'��K�P�mo]/�H��Q��T�&㙒�{�j��a�i��/��C�ٜ�%"�ĸJ��j���4�����`�Е2���I����-��0`ҁ�6�lbpY���S^��Y�a.�2�];�dƃZ�d����º���X~����r���E+C,�J���#p���FG�+G�Y��=���[k��?J�[Q|�ex�J#�[^��GþJZ�$�8aE3!&�N�r�X�C�e�0s�8Xj�PM����~��B�q���YmX[A�2�IF@�ym.����K<8��c���L"C��_�Z�.���5�w��5���((B�Dm�����5��I����e�5ʙѵ�ȿ3�Ǣ��*���������n\��G�ڣ�.o�����b�`%�o��|�fY}kצ7g��T�m�4s���rcU�>�ʱ�p{�?{���E��BM��'��1�l'������rƨ���	I
�; `8��"~�XM�*4)�\�� ������*`��7E��O�n��S��=6��+R����s����C�O�.iw;
���"+�67�#�"E
.�AtvP*l;S0ȵ�`�Ik��[.{K�f��?�O/vs����鰬�3b���q:����Ғ�58�ER�gD�K�o�&��:y��+�[��mٿ��F��A
ĺ�2`�(7di�6p8#���g���e��DS����p]L�HK#(|8KI���/d���d�e�@c@�ݳ�dcD�y�q{�i�����"�)�G����5f�M�Ԡ�.�(͖�i����1�q�U��keQ%��uF}�6���t4`7Iw�
�5
S�Ök��cxʫ��~�����N��yk�E�h������rغW#C$��._����v�''��
x%c���ϼT��B��w��`O����}>	LA��Z�[bE��f῁}
�;�/�� �u'*�[c�fU*��K|�׭��� KН�F�nn�Zd9��������H�
u��O�rr����A'��ޏFOm�ʦ5�Ze�A�^���9T���Q�yYQ�2���B�\}fS&c~.:���ݜ�9�ᄗ�B����;�B -��rk��_�ņ��^�"�T>f��}`�&i��a�jA�j>$�ҫ[h }��+�"����_���V��{]�ˆ�ϑ^ո�)�+!����4�
\dd�K�B��3R�y_�����~�c�a��i��!8dy�f!�$��6��ܐ�|;���9ϓo��{UK鴵�+E���¾�|�F�O�%��:�*�#�Y$�ԯA!�w؇����4��wh�i���̄an�s����s�+��Y�d���K�R���0��_�#ٮ�B�(K;v�b��5~9&"1�z��K� �qO���,N��7��"T�4],��08Z�^�j�r�+�A_�e ��Q���*������*M�X�)O~�L7�I�lHQe\ �D��s����ƾ�0�ۗm�
b`e���ΤTu�\����g�:��R\�jՍ�����C`R�-Zg�X	���b(4��W(zQ�3tR4h�����ښ ��A���Sw���	%ᵕ�
�����Dsp��J�%����eh�	X��cW/v^iA��(uE�]����eli�S}�q��־~��}ڇצ���E0i�'n�y%Xۂj���A�.P�dqFbf�g8і0��3gb�|�q�Vt^l��
�fl׼uHd٢ ��c&@E�>^��w��q�䱆0e*�:�uUg��P�l��znE;�l�5~x��!��q�oל��C�A4f����ZY%�˜+Ŷ?��_:��,U�����|T�e��l"�h7���7Q�
��wϰ9���J0��e��3��#�hXgb!�qځU�u�˹TG�743��7�y�j��ĝwkh�{h�hP��w	JG�w���ֿ�i��Bt3��U���J��h]
�Uw�p��L}"Lr*v�I��������8wwF�B��/�4��Q��5Aw~�l#װ���m����&tM�}Vx�"�&|�ʶ(G�mz�/�U��G�;��xn�U�`��������| .��E��2�v�Q�Ӫ��@����͛�8R4{/��#<�-��U����r��`ԉ���a��qa�9Yh�� 5�����D�&�ˀ��^�pϩ$t������1�r�؃��M�,��=a�zѕ���e�z�-�,��e�G'^V�)�z4���i5k�X/��=k�-L�qC�����+X�@�k��9�� ����j��
�n��[5x>�ȩ����u�O)[ȝi��5��t>�׮����!l����[j]'VC6��K��~&�U9���P.��~���%#�;�}I�-���^�8v���7�_
��i��\O1��2X�2*����y�T�th ���x��F�U�������^�I{ /Wϲ�J��'_W��W-v���U�_4�ʃx���*x?i�� ���}�(.�n<E_���3��'�re�14Fdm���i���Ny�0�]w;�d��+t���]-�]��7��Pe�9�I��E
55�-F�Q�p�!�q?�f��6u/7�InG����.���!�h	����~U���q0���?��vV����M�a�~���$Y�h�ݭpEsP�\�?�ρ�CH¦r���Wc�ҥF#qe ��`�2᛹,6��t2ߋ���)�bK��Yف�(�����uk�.����S{���B��,9�H,:A��S���_�-���_9V�a�=R�6����D3���ff�_��ϧp�6!Ȱ!.���ޯ��������:���i:SM!��(5<�S��I����[љ����Gv�:3�\�+d�Tz�7s�m��	�w�i��Y����{��)���\�K��� �
*�o��]΅�r
W"�����!�9f\�����O�GCE�
lR��؛�/���$I6x��y$��M�9�P<��z���ွ�L�4�GRL�q�T�������:= Nݖn�,/KdX��OL��L�O�Nx,C������G��
�:����R���{*V+�2=���W�ҳ8r/�yHΩ��mnNd.�]���"���W	��� 5>d��b0��*Z�DAsu]�TT|ǃ�]��K9	����!�-ﾨ��fe�֚��'�t�c���t	6����\YG���as*�����c��y�à�.had127΅��T��R�	ķ�P	_���e�%�E�Vn<z��1�M1�ؼ��=��5D��@7�H��(7�⶘N!�!���q[���_UȰ���q�<�>qD1@\��EW� 巫��j�%ݧ_���� �K�Z�A��͖�V�u�+�mRA��^�0/5	J��/;L`9}Y����8��@���%U�z�@1��� �I�s�#�w@v���ƓP"+_ପ�Xr�{�ʚ7���!8�{D��e'v!z�XI���lJ�+��/o�zc�$<�x��������=�9Ah�O����u��OK2�;��C4�i��~-Tr�Kw0[8���fO'�o J������F A+2�������Т�"z=����T0i���&��+
=}�!��vp�CO2���nኧ݄ TK��Œ<��tb�]k�����`V���]:�;��7�
\���٘'s%�����Z��3���_m�E�F� c��4�qy<����@A�>�Ճ��$��j�iF1V7d��,Rx�����`�B�@�
A��2XHQ�/v����d��F�P\�h�^�0��z�Uȧ%D{��'m���������MoGR�!�ɯ��5Bb /\CPk��v�9%�� ���7=%Q���
z���
}�@%ph��j��$����IץC^�.�=Ca��X�ؙ�q=]�I���q��Չ|\��D���J�7�1O���S4��[��i.d���Aa)�p�f�YR�t��?d���`S��=�����G�?Y�%@�i���A�˖b����t��֮��o��e$�5�>	g�F�,��)��VF�&яC���uP��������6/=�E�d�h�|��� ��]�d���I\ ��_1ޓՒ"�[�Wrw/B����cE��Go���ϩ��J��M��WŚ�8��4�2{5$M�F�~�<�uWJx����ܻz��JM7o�s����'!}R`����g�}X��i�gәLf����@ݍ!B̆)"�E��K�p02��P�u����+Sä
�3�:��u�Q��?� �$����_���w��뤇BS=ϗa�.h#�{a}=�b]�@�%�������!���"����g�o�Ÿ����8�:��r�"��Y.�6��p�c��	e��S}�ҏ��m����6�ﮥD�F��V��\�5��^�ɓ�ǘ�#;��y���]'^�~��n�yM�e^9�R�����A��=�q���e�����z"m�^xvv�*�sV��tl��򧸂HݲLOzs.�%�
 [c5$@G���`�x�	q��q�Q�d���6~/iP��g���nyF��gh�hѨ'&�|:�,�9z4D4Q��S�������Q����-B�3�������U�\+�R����XZv��Z�U��jS�C�
K9萅~.�����^��0�D��H{��c���y��+���1I%���q���sfc���:��r���l��g�!_��C�w[�*ٴ_D6����`���q�ӡ���6����$�M�(N�� ����v/󮯇^𔖗
rǪU5��'������������L��tUg��O����T����m�r���`��T��2D\
ѝ�f+�'�>��x������X�%�	؋tNKE��p�]��V���(KK=d��uT���"����c_҇�0�������֪�Z��5�2�D1�qB�-�g��d��1��'z�"���<PI�4�@�!l�"����'���79�`�-�tY�$K��p�]'����k������[msn�P�T+��c/��s��sR4d�oq^=�9��šLV�b������|�B�H�����jf�S#Q��M�ZQ��P%I,��մ	���d~�ݬb���l�\�&�ݯ5�a�ӗ����.%䊶go0Qm?����B�U��t|�ٲ�ףjS.��x=b	p_����V�7�,N�љ~Dm�	K�1]5رSl�7|��:�Ι�эkB$�}|�V�n��`?2�R�ؚ
6|�NK|MZPv 
�E�%~�l[�đu�tھ�5�-&(�:ɨsR�ʁ�g����A��7��y4�(\:c�h�GB��^�ʎ3��Fa�c����@�
4��kF.'���~�#/0Y�b���狭����}���
��aقy�E����1Ƨ�M��^��\
���M*Rj�w�����*�3k�ʂի�**����]g���˜p��"�:M�筣YRYaDE��l`�x
<�eԂD�����=v6;�$�J��m���IP;� jS&(��K��v���Gv���'������1{ɜR2�Z&�6^�/d�^����|[���ewA��t��Ibى��q��%{��j@ �]�X����u���N��Sv�N��,f���7��*^�ЬD����ʺV���{%��̘�[G��yMm���d���{4n�n�n����Կ��к�S���+�.�i�9����*�;Pܲ���ijN�~dې`�W2�	>����
>(�2	ء��c�^�[#غ�g��.�@?��t�M"D�\���"������1UE��q� ���IJ�\?g��a�h䭸��Rx$aR?҉��9���V+�db޼#pb��%5�w�h�`BJ
]�=�Y�"�|4�u�8�vϴwp��I�����8��5m�ϲp*�Q(X�hfcJ�yXH��d�:��	B[8V�$������[��E�O����Ȅ�����v=�o�R���R.fr�Ѥ1�Udf2���pP�&u�-��CÍۋJ���1�`��g��h&z$�bV�fݑ�6<���>�ބ��tЈ�2�i���a�;��w���f��RP�b��;f��y����E��&y<4��/��~Q����7���yH20QY��"��K�C���esB:}�
��kҟc���+�?c��rF�c�q0L�ڜg@p�TV���|.��:aw���ԉ\W5VdX(�B��]#�~C��l��Ulk���� Te�.�K�k�,�rL;R�mi�� Ғ�� �C�JRF�V�����;���3x�Eh���թ�=,��y�� ��?��G}���Gy����������bi� P�}������"�=�D\aL���w��{���Yūgi�;�jZ��蘝��Xk/f��	WrӪ��'/����`L����(�yavO2U�E����bdn�	��?���69��0622�.�I�=���q�FpB�<ﺣTy��K|^y���*ε�����
�r
+9�
�	��#��I�XY�F�����ۗ��Z$�����-�Ÿ4�c��َ6X<�1�0[r���P�ܭ���`�'i?�t�I>�@�b�,g�oU	&gq���"F�>҇��0w�L�x3��%lU�v-�t�h��/�+h�$���>�ϵĝП�r�ZU�>�x���r�6o�A�w�*Y,��D�4��@Ou����wH��8�s�u��)�)\B����&��Aa}\�Z��8;`Q��I]K�7�����@5�m��N�雏���(���h*�o�"�ϺĔ��2�+p�! � fƟ��%�.#�������sZ5�6��,���')��a�Z����xr�;��+6%����1l���` Bm�C[t:Jʋ�
�s�U飂c��]����\D4*�S��k��?����`�A�]�S�4�Q�2�Ⰸ��;mҞ��T� ��$�=������A�ɵ��(wuw�X�l����+�ְ��;�H-���j3�s$7:ZA}X�ŃHg�W����kڟ�8A	�]��i��^��B1"�S��ٽ ���ݘz�<���x
�
�>�֊z���6��c>���l��즔��a��f�|$ʦ��MċX�5g}.�AC���x�h2j�-�}�����)x�Ô���D,���KxY{����_�a��j���=�?É [�A>��q�!ڵL������\�g�-3f������Ҧl�@P7�T��xo�k����Ε4{X ^����#|�jknz/x��� ɕI�~=�����bRޚ�7��'���	��\�],'��W���Uf��>yF����A���ן�y��;��&���f5�Ũ]/�Ǵ���t�D��K!�2�Gϱ���^gyN$�*�i�yy-��Wa��]I�`���t�U����D��S��;�C��%�@1��/,�3�\�Dq�S �Ʃ'�(��	N[}���\�0�ӤsR�*T�5#$�b�i~R-
�4��z܃�A`��-���*3��'~3b�=�s�LۏĘ�ӊĴ->]x�9���al�ʀ�: G2^=�Y���m4��������Ƹ~���=��� ��|n�LWZ�t�J���<rU��a,�z��q��U���B�?LjЇ ��+�X[�:�d� �� ˡ]R+;��c3	�+c�����.�h̓
�{4���H_8A�-�+�� a�=[��G.XՌ@V���0�TR�x����8I��8�D������CG�8�'ҧT� �rPx-��μQ��c+�yY�����T���|?�����(%��˞`�m�2�qI7w��T^����t�ݶ���m��$���-�KLt�]�.��� �;e������ր�Awc��i@�l���9��?I���T��p�$z�-M�Q��;O�pp��w������,d�/������Z@�&�p9��7^�wUr\�F�V�2�Q��)�.L~Ƙ:DӾ4�+�25�?�W�A�xƎ1��R�{(`֎���~�����z��
$]�G�.��0��~�}��t�i�a��II���pfhnׁXRb�.�#YA��	��pQл�M�*֩`y,����S��Ӯ_�� ��Ǖ�ħ�:�rpt����c������{����@���вf�s�u��Ďa�8 A+@�����H/�� �q�v��z~]ީ��g2�(��P6���3:��v/��g���w��q�Q��(_	�.�J�� � H��F�y�,'��4�S;nf�ȳ��O��֬h�d�07F9�;�@l@�&ߡ���<�d�D��9�;�Ѱ�eϪ~]��#�cZ��{ұ�?�;�-�/�� ����|l�;���x�������U��H������1��6=o�-�$T�
Q����0� ����^��'P�RJt����MS!�P���hf � ]����of������}E��c"`T��P��������Iǀz cpŏ'W�3J?v�W�Wz��2ik�4�k���f(eMY=���#S8�ED�
b# �`��iI-��,8d�niDz�j�;�6��%+\aP@8�	�`���b����K�+R�o"����\�UU��X��hM0	�@O�����t��P���}+\�K�WO��hUaRnS�&1<h���*8N}N��"�ϋJ�&���C�Z ���M+��:�U��%��_��� ��R�-���$~U��H)��0�u]�hx�����ؓ}�[�ψ�����@�zT�iTz8�m�xsg���i��}�ՌW4~�߹����"�;
qq��VCL�P$go�����X&>��b���YxkN�Ђ74Y���.�L�TO7��>ߓIu,��<E�ܚ���yG9�0b���C�U�_�	������\�!bϽ�ʄ�Iun��YG�Ò��B����M�����ה�B8��r�ε���Tf9������9��yB�V�lht��T*�ٷe�\���n�.�� ij��`���%�d�X���~m��%i�4�|(jn3�d�yo[Jj�J�M��������N|�︬�N}���Q*l�O�@�ƪ����5��>gg��Rz���[� /n����?>��+���Ez"l]ם�:Q:�\�)�J������	H�lU$.��r���NA�\:���0C�j,h������54��j< ���/�9u�",o
�K�FxI�_�94�]�K��#�E�>@,�m	Z4QƬV�	>��G���'Z>�
��ڣ�2�O�Z8�+e�����jr������1�$!#gC���y��\G��B��09�[-5�G�I��K2,�ӑ ^<�^[5{%������_?�� ��ZIܱ|o���%�\�V	E�F�aN���p�{GS$n@	
��[@�TKE��%%�#S��p��()����I�~@ꐲ���a���͓���i/ʜ���0��A^����D��ۥ.�99�#��G�tt (Ө��#$��e�P~өx
�x��*��S��ߺ�QpF�fx�@�z��G&;�����X:���W��.��)J�SՈi�#���ӥ?QV��*R�FB��+��%O�BEC�5�81�L;*�������.�U=�p(��i�9+I�.	~PL4k�(�+0��Bp���br�À5A[F��b6,��Y3�4�щ΍��,\���heC�����ߧ=Lk*7�P�"�H��q�8^���"�R�&h�P� ��U�E�^�>�F���M���r3�CϞ�&X HA`���?��W���k���l�?w�)��߅��SO� ]�g�~�N��<� �%�iI�z��TA�G�MZ�,��rEb[�'�x���v&Ѐ�tR@�ЙӼ�	��k��
PV�|N�y��	 ����߅�V���p���L!��b]��s-"�歬��~]��f]K�a�ib��[1c	��#F���PW��'n�G��4'����	g�-(�ݔ�v�p2������pD���t�����_t`�>4�� �	��c�����(��D���-0+Jo&E�T� F���^Ň���MÌ-�B_�¥��Ex�1���7�'q�����ϱ;���!d��oFQ�?4�9����#��~��U0T\�㏈-�$�ɺ�wR���!�	W�F̥/F��v��NU�J)�A���Rl�T���E�7���Xݥ�=�վڀ���M1C�8��LƵ�U >���y��+�̊-=@+飲ĘlTό��Ա<K=�M� �*�З�.�F>�Gl�9����b��.g.=��κ����7�*ܛ�f�z�U�ZE4'��F�Z)�*�*�؊�T�H^�s�8����P�j��(u���s�4�}}/����氾k�{�߃?��b��p��	��^ah�+x����~�z��<p�2�����%)f�D���C���?MB�������~��Yf�V��J�W$��K��v��Q6n�K�f\6�
g?�z�!��_�Ts���:{c In�t6���Ne��ݐ��˾>����Fg豻~��+����rQ\�*��~ht�%1ŗ#���K\��`��r���s�c�u#J=��s�m6mM�͚��&j��0"#KXI�MaB�g��Zn��8apɱ��[�b�>�Ui�C����/K���SM�H�߀3���T�c;;��G���Fw��P��񃖩����(^4^ig��˟��faC��@�XH�}�69QAe
�ҧ-�l�҅��[�A�nO���˷�h3��I�n��e1��WюN��Ü	�LT�,�FM�:�s��jR���r��1���}J�P�~sי? ui?>H���\�ǽϢ�&�XMw�+P�Ti}��?���ڐW|Y�L��/G-�� �`��!��62���H�
oK��Ө���c�>�F��ʁA���md��Fʯ�@�5O�=���R��|��$&��ю���d�.`�@X���e�q�2A�	�;9��ص�ْ�@��7k{��mH�_��F��TQ�UZ�-,�}�o?�̼琨�^�r�2�`z���(�`<�lJ'��z!�����*ǁ�˱�_뺙:��^��m-�j�J��̨I�5�]���r�pN�Y�l.ڜ��=+_���;�M�:�ş�G�=��!�)u\�[pˋ��@e�*�LUU6�\��r����&��v�ɍp;��f��@��|��#v���-�ww�e��č#�Z��W�f��U�";��"cbu�������&FZTՄ� 5A�<܊�"��f3}����C�=R.��T8�z7�?��L����
�*H���ٓ��Z�ogk���׆��ӻ}��Q�*�!*�P!,���Tj��a9�����{Խ���{��O�_A(����?�(e��=����I
E��}�ztiA��	��@j	�vpI#P@���\�Is����S���`"@ȜNX"�Ǆ����w�g���sS��Logn�ƚq��]���؎X;���︪b�����2]14�]�����	� �g�&D:��My1�G�y#-��� ��}���1J.e=e`�\v�H�r%��/!��P�q�x�A�_	N�9j��xkR�/?P�U`�= �o��V��^=(ttvz�o��n��u�ehg�Zq�>|ނvܔ Y�	tM\1��i��L���*��ulG��bs���檫���밣B�GM8�E;U�����(��@D�8��57
:��<�.p�7�����Z>T�q�m�mB�j�R�����	�׸-�Kh�L1;���Yl���FRk6���4_���R7��� f,��U�\
b��F���U���Ӱ��s	�{���A����!�B�0f^6�Bn8���on"a��E*dg+��هy��owؾ�ˈ�p���$�_�/&&מ��3Y�ڳ-�	��f^H���$�u��{m\�B�_���� ���yO��n�LՄs��Њ~�剂��ߠ�Z-|�!���S�X����m~C��Z��݀	����{�&7����2C��Ly�P>��bh��i�O\����䳁h���vCS�!���5������P����Hi�=�Tݷ��h��!��4�t���I�`���M� X�[y�Q��^�O Kc<�ӆ�
w�� ڬu��Os,���t6���V�/�uV��+��~h��YI>Qe�:V||!G��^�Esr�'���f�wG7E�O����	2��ς0�ϡmO.�~��&蚘���-1�[��q��|-bӊ����޾Sʴ93\���X��	�����c�m0�[d� 0��E.�{`�h>�X��o���"T��\��@9�8��2��2��l0�^���:�o�r�h�P���Y�Fm}�oo�M��+�	D�86�.n!;zdw��K4a7�,8W�!0z!V0���8�3�%��� u���i}SB�I�@�J�g^�(��^P9�Ե�������Q�F����,�������Ki�-��������?�>�0}[�sI�Xe�	��~$�m��9&zPZ)�4Qs4�,N�>�튰\���:<��Z�A.�WmRa3)�n�[�%�0l���rz�5�~�B�C&K���R9�Z���.Ĕ8�#GŹJ����ݖ�7�m_/\I�{�Бw �ݬ��301�|6:!x
9]^r��OU�/[A�71+�X�CKu�̧*~��u7��j��lv�$	��t�wX8V��P$���O���նA��D���Vqm-��LN#�j�	��|���� � o�lO˔�C��F�})����5�U��di���j��m�Z�>4;*�zEߚ��D���%��I~PeΏ�b��\�������K��������4���9	��=�M.�p��6L�5ų�c&�`7��O�U�  ��+�]�;�șm5�f]���7��q0�C���o�pUYŶ�:�&ʺ8�&�?[���1
�#B7e�YV�?�q��u��ۀh�;�b�Z�� P`ZԎ�.�����lF�3"L��e�,�t����4)��P��-�Rc�����R�v�)M}��3�=��n��3��Y����-]��N��?me�k��xr+��sL._��jF��,�s[n��9�a�o�T"@������Ȋm��a<��4�^�җ!�D\�o��9�{N���1tp��D�k,|-�*��-�R�m�y:��'S^k���ce���S8�LB6�5��("���f�%Å=�7����~O�Q_��U��rqyy������I�f!��7�������{�Q �Na㔗��{E�ᨱ�iL�����F�3ۥ�fW������ن�����vz�^��U�9���y�W2��4\}~�B���h.l�I��]%C%7z�5��^&q���Q�mu�q��غ}`آqă�T��L�v@g��[ћ�0�]9�~_ʤ��R��
l��X!�t?�[(]�j����t=r����!��ٙ�[^͵�_Mk�;�׼T� ܿn��8�/@e�(�*�v���;oD�.�p]o	�V�#��v���S����3m9bqp�!�墪s'&�,�p������l����6�
���>��M�/5�=Gni�"���DX��{PFy�&��Z������y��+h��C���d��������*.�)"��L��5���;)%/O�¯^?J�oh�b#B�����kVw%��O�Ő���R��d˔d�Gse�^�����~�L�#T,��(�J(�O�Bz�z�i���".* ��5�3܂4����Q(�&�"�D2
g�������������O��Uu{cͯ�[�ء++��+
��4�a
����a�8
z<�9�?Ӣ�F�ϋ�R��Ap��o�cZY��D��h���=Xpx��l3����.�ψNV�*iZaݻ޳�Ͱ�ڣ�K^�3��������-��B8&��u?QѨ��x_銌D�^�)�;Z�SNB{�����0�E7j�0M|9pl��]S�d?4Z�n�a=VB�T�Q��D��Cr�@�P��2@2�͑2�\^(��}��x' .)�(�GT�1/WVI�)Ur)�V����{k
T�
^���rՐ�x�X��<<���}d��݆�����仆����=/��"��D�;��ys:�<y�SelX�z�tQcϊȧ�2;�^`LG��kH��9�z����2\,M���dk4����[��T�F����	:ۢ���CgӞs�ֹ�)��7�*���z�bN�_��6���.4�6�`jg6u����˪x�9���ս&?��������r���D=��qm�-2�h���2M V��t*������6�a���3�O3���I�v���H���\)j{'��웥�!Z��4�N0�0-�[vbЭק��:i%�I�1:���IN��폭ʆ-"�ŋ_D �*��a��������J90���IW��2���^	��*�Du�\]T�\�g�3.�	��}���X�q���b9ʺ�U�w:a$����C����и�	ǉ�7��EhU.��7�{|��J�������_�+g9u��E�Ki��z�,�N�A�����BI>!�ᒌ��C��`��m��4�2�s_�8[�Vx�!}�c<��>�w_|��O���K�z[��O�?�Q���HQ<\�%�H���ܐ��H�Hg9�����pʓ"���pU=��������V�<�^�������ζ��l+`#uMX0����|(,9Dk�{�LH]����G���q���|�U��P�-�A?�vᜈE��?5эN��!�f/TF���x�+����0�� �� ��`U?��%�v�Dn�� �^n^��z�P�
)l����53�����slNq���XهO�5k�~��8+u�Ƃ׫n��g܁FI���-��6׽��~v�:=�
ތ�08t��EīO@[��!=*�o+6�aͯG� 8��_�9<S���$+~�^.?�s��G�t��cKA�%��"�[�H� ��ѱ��DH^��\���h��š`DS��S.?�JO8F�^^{/�*���4��+2+�5�;�h�k$ei��D����h��mr^E�#QW��C�7{�8�,��q�9$�,L�`�6�嵳{�2��ɰX��ۡ�DgJ?T��d�?#q��"}��V�3: (o�F*l
Y���X�9HZ�	�G���>�yi\���`LZ��:�9X�������]#�P�}š)��q��U9<��U=���'D�[�����}(ʄ�^�ף�������K𱏧�1q�R�'���i8{	'R�q�`��^I�ِ_�\;���Փ�j� \���V��#2I��-�"]<���YG/w[���Zϑs�?J���
�� ���0��M����(4��$ P�K�*�DT-u_酊�ܦ؊ybJ����<�Ez���@A�.�&��\�)5�h�������ڍ� r����rձ��`�ܷ%����E��^{������}��6���%�f$i�w�`m&����;����=t�i�pb�,��-0�����6��h��};Ի�Vd��b���bl�#UW�;��k>D�[;�.A9:]��yd��̵�gh���/t0��^��}�t�-��7vd���y��DU]m�yH4r�'�3��f�@���/{������"��瓑��zἻ�R���ή��R('u`$bQ�u$�X�+����L�����|�-�v�Y��oI+�ŎSޮpݏ�,&�^E�E:�A��08�H��-C�g�}x8��p���Y���E2a�>~�Z��&n�P�I��FJ3��I�{��N~]=-
���mH�E7r<{��wA���la@��=P���?!��w90�͕�f1>%U *<����y��lz����6ǉ�Q.���P��)ƕH�*��`�X�n�e�+��ٌ�D�q�	��"U��BQ�	�ZH�����Gg�aZ�[�o*�_���+]�����(o7 ���}}n{l�RmڰX���5�w޷�#q�0iN/$juqG�x���a����a����m����5e�ͪg��|�|��$�~g��zh����K���J^�h�O�~s4�6�h�*������Rq �٨��E�9ӵC�&�Z�_GL��K�������v�{�6�A�i�!���%�Y�0���*�`�k�jb���B�+��(2����Ƶ�2�859y�7�3R�A�9R5S�c�!�h;�����d+�k؂u��9�rxZhY�(a9]�����9���N�W*���M�����Y�2�>��0[`�uI�ʤWYk�eٖ$��J���@���@��O@6t�Y�ΐ�'2W@AbY�H5�J���Ƀ^�ꞿ86y17��%�T��|��r�4��Ql����>�px�b~6k ~���[7����rR)hu��6�P^�r˪��JR��[�e���aq�
���0jZ�=�������۞�jmƼz��8�RW?O�`��혉��opn��^t*�W�ۜ���h�����Q�v[Z���ѹ1��a�2'&���v]A�'Yℿ�I�ΦlM41��!�ookBQ�á}z�«�5�	�j�t������JXA��9:t�߁͋�3J׳���F�LmN����aQ�L �S�3�e��L�4uQ�u�w�������0���(���h˴ב��� m��v0E��D������4���]�z��i��{��T٘�J����b���G��k]Y��Q	�+�y�*�Z�n���Qta�/Qe��!�T��|���*:7�1Я�J�mf:��{�ʀh�?�#tĞ)T��}/��\����*�|M˟KC,mo�ޕ��'�1G��R�ժ���d�>@����F��Gq��A�q������G���&�O�n����G��~��^�Lg���e�=�����e����x���R+G�Q���<���讍���i�Ɓ��J��Ft�N1b澀T�����(�����叾�a��+*`��kfC�U;p�Z-9Q��1[��M\�PLZwe��zňKji'�R���z$��R���P�]V}q������Z��%�Ƹ:6���Z�̎�v<��%E#�ư�j��
IӐ�L��a��I��q?��p�K���k�V��.�Rlf�������Y���[u˘f�)���f3p��/G��m.rYV�+�"^�/A5DH>>=#i�`��Xb:��2���){���p6}����7Q�X ����woWe�L^9�8��|X��c�Cr
�x���Q&!xC�N�)��I{��̅h\ `x���~Rz�:��O�Xo�˽�*�}�[�D�̻Anc��<��+�h��J�"Gmj<�X��?֌wv����x��y�A\��?S���13�C��8���ċ�~�bts;Ȧ�Y�Y��9�f�]����Ͷ�d�����K�|�����;����e��}jh��rW����F�h�f�d�O�ߖ��t�#����4�:>?0����En4��d�\�q1�1�8���V��E@ؿ�ۇ�=��?K�^;��ӽliZZV�HD[����W�!7r���X��Y�V��o��[�ua�@{�2b���9ԷJc��Co�����\X�'�t��e�@k1ԯ�b`D����K�m���2=�#�JRL�W4�4�x�+ɜ�������������	6��_����� ҍ�y �U��tữ��316z!��p�rt�ŕ EW��;S«5����
�7s�(���}��#	]�+�r���h�Y��C��vE	�c�c��Q!Hz�_� �X��>"�M�=S��T���J�o�M������ѹ�Ea�Wy=��.�}n�H���.sfoR�	�)R!�w/����W0;T�"��^^��wVV����3�^��s�������&ita�Ϸ���2%�����Qq'K��2��s�!��7�q����_-��$����[��'1E6�F���5�I���� udǉ��4Rm�K���>��6�_��R�!��iOY�X�S~ǿf������Ym汑	w��Y>u�t��1�H{z���x�6L�xsC�Zy�0�-gt\0�1Ε.wX]|���~|�#�:��"�e< ��A��uLw����G�_�
c欥f��+��}�o���8��~��	�0؃0fAv
~�o�]�����}��G�Q��/�vs�k<��YV>�_�G^>sö*�T#���4�����.�1}�2��Ǡ�?|l^H�>� �｜[;��|QY��ڋՊ����Axy�� �fO��g����ן�R6�A��<�F) �|�}Cb���&䖶�,B�w��0�/x:i�C���_p�8L������d����u�KE4�}�=eVPA��G˴@��wtIN��g�Q�V����	�G�V��:%�M�r��85��y���q�}��K&p���I��V�_�1U�}2�H�����R�9\�~�_~�mƆvդ:������Oͫmen�	ڠY��>�M� ��^y�$����M]q�U��Ꙏ����� �ݔ-���E��t�l���n��NZ�`�N����Ȳ� H����i���c��\�C
5�1��o6��A���cg@ Vܕ����b�t���0��Q�/��k�r�,�����,`"���ҖvM���v�WzșX�q��8�\m�Ƀ�#fC�y(�u�I��h.� z��B������+\�a#�s{�'��r��c'�����K�2�jK�N��ق\0'
����[ĥ�~���۽���d-�c����M*Qk�z*�%�@iZQ=�2g_���0zNS�ҳ1����k�w��T�p�/L�������N�e�3�_Gc�����	�&��7��Ct��Ig�X�$�u8z���f��|��CP�pOh�E��SAre�;��6_�E�|�Y���P���I��fH��^D���j�ҋƭ��(��R��Q7���
4-�j0L�����{�����;�]u��$F�����O���P��N�!Ki�
o#��r���g�މ�:��wC ܲ���,* �o��˩k��m�KM���s��yl9fMZ��}Ą�ƂLE�8��Na�l�ժҜlڈ9Y2��9��JV���B��KO�&yC���	5qa��0��l���o*���*;r#?>���JdEYV�<��|�X �R���<��`�
���q����Dr@X�m�i���Cѯ��|����Ŀ��Vy��pV1{0ewV��]Ll򂤔���5Y�N�C[(z�9bD��`�ᅈ�?FLy���e'!���3�I4�K��`H3M�9_g�垐��Q��ٓNǯ<��+�	 ��:`�C�6Y�:7B2�[�J�� ��+=GJo�P���U���>�n4I9Ii�c�dl��
�fn�]�O�[.e�B�r�ϳ�$�������,��)�T���y��0�y�	^y����rY[t�iT	B��zQ��������H�y�n`x�@@�9�^��k���!�� 2�g���u���XA���ڑj~Bw97gB���I�#��1�*7�\�d���J,�*:�K�
pk�>=0��(yZ�}5��� ʇ�h0D���e����}��^'io#آ���H���Md���<�ʸUyW�Ǿ��۟|
\5(��f���7�|ѽn�&�m���ro,S.�V5�|�Ӥy�.:G�|=�)���4�Qa����A���[�Y��M3�O�E��ʺG�S� s�7��0��NL��:'x��Ur:mHR5>��J2��h�/
m+��?�2����R���-o�h�M�ށ?0�e����8��=i��i�q�[�����.6���P}��Оy����X��Pٕ�8I�[@��J���[u�,Sy ����	�1��SU�����x�Űa���8f,�UW������W&Z?�{�f�\��:��om���[�7�GD�D�<�Yȇ{}TuP����� RE22�?#G��xߜ����N|z�7����}�p���/p�H14z�L�_��'uϠ%!��a�Ͻr�R��Ho�sܟ�E�Vr݀��֨��5JnFʖ�sU�0~��:�KL{6d�j���#|��|�T��:��5�α#���7�I���]�s����t^q�A�h�Aɒ�>����̍� U�Q��L�܊�	X�Z�q �v�����o� �G@Id�|�^q����z�'�-���L���0�2i�ِ:��r��+�8=�	���F��*Qp�O3W~te�<C��A|ؽ�i������xB�C�f����v��7;�
��<y&�klӆ� I�؏��mWG�UmtC�FM�1[����f~���e���s1n;$P�����_.�]|'��{�{�J��KLf� kNm/:��3"O��`nQ[��5�#���]���9��i���� �����G\������!j�'����_�@-;ǁ$�_萴���Pf�kȻ��T�H���Ü>��uL�y�ȁ�r��X��z@��~b���bw#�D? ۔�%ӌR�ӭ'N1j#�� �)�&�&��]���A��VA@t|a��7��G��!�]�5�*�Kf���H�]�0B�[𨨬��^o��I*.]w��OI��!������P���ə���I{��	���M�� ���odš��wZx%�l�渷�cr���r��LV��� �X�@��
���$�u�#{��#Sφ�uh�z'ZO�:*eU�G�/|ۑ-f2i���Y ��̲q*��)<��u{�o[���J~�`E5�a�DR_sg�����O~�˕z~O?$3ͨ��[�.1���`�F��o��̒輿��F� ؄d�r����y��(�S�������$�g�Ut
�<����<�9�O��������J��Ď*ft��%��f�M���D���{�z 9���v\t��a�9����?�[U�7��eNc�K�z�?~�5�V/�����:�J:8��Opa�+�P�pH�_�3�l\ʨ3�0��P�f���͝����Q�0 �0?�F����,
�<~��-�l����۝������0`^Z�L�Bgl�7ȏ�����N��[��_S^�V�>6�����	�_��h�x�m�+��(�.Ik6���q�)˰���⟲��e�&^��M�n�6Պ�]-{+0���&!�z�.G�e��j��'ĳn�?�8v�LÞ�����4�M9G���#O~W�eR�v~�q1�\��p�*�{.ck�C�}Q�bq>N@0��<H���27�	��h�}��ŕ�t�b]Q7��&+��Fys�oS+�*�D��B�s�+��r�Y�F�L^։�)â���@o���5e�b���G-P"lC���(ǣ��K4~��V����Z���E-��y��%r��gC*}MC���\0 ίDkb�gr!?{�I�k�
$�xK�/D}�I���C�8>��U/ER�8$�QeFW��!�������ą��:����&w_\�i����mV�IE�iV�F0]+��[�A���G�,�}������e=0���N8�4��6 ^@6�$�f)�-�_v�8a\Z�~JP��Twd9\���(��U��S�,�A�����8*��U��������W��t���E/
WK�,N���R�d�b�2�mE7Ͱ�l���|�B���i�l�	`� J�T<R��~���,�����E��,$�\~F檺~�Ű%)[�(@^l��<N/����@���Ht`f�]A�^�CX��8LY�Z���W�k12bح��3*F�MnTh����I�=c�n�G����{�-w��3�ᲇ��kI��c�W�D:�ݧ�;�8���_�~�!���T�2�Zpk�n��-��8a���8�ɔ��0�!�Z����-K�6�9:�����6���W�5���L祉��/w�q��7��*Fx�M��l׍<�*�=�v����Έb�9�ܛ��o��#�RuV�~Rvc'>�e9/��d�CH�w�Lz7�KS�G���f��g���Ú�ڌG��-?�2M�t
L�p >ܢs~����5��="b�\�e�X`�q����R��>3B����l,H���	�q��.�j#$�5�~��z�2�xR^�$�ͩ�[�x���:��u|�Յ�� �����	f^l,�i�x�D������oneF+�Ł��Y�z��
~���jXO�3����ށ�r��%*l������~��ظO�D�EQ�F�}q/�»��"}�Ҧ~R$_Mk��o�B8��l�徤wU�z��,���&�<	w�@D۪�J�Q���#���8���Gn�x�R��80��y�G3�6��4�/������1�]��~I��X��҇s�;ؙs���:������>��x�[�W�%��f��SYz���|l�F��H�1h���3������)<g���L�-�����'(�� ����ǹ���0t������s1}�N�[��&�#�0+�!��Ve�YR��\a�q�ta��FH~���2�<�n98�^�!H��Ũó��;w?T"���n8�,�:�tT�m[c��c��bݹ�򇗈�
��忽I/� �%X"$����&n���ҿ����XJ��]�E�Xm�6�5�LO�ԡ����lѨ�85��Ǡ�
|��@�qR_�:8Jv�XVh-y}H,�]��Kj�K_�P��KS��4�[f�5C]�ߙ[���%������ѵ*�|���U����xhC�Z�zk[��^r���w^֣�΅Yp�JW����`g`o���yz0��|[�3���
;�:KP�`w�*�v:�喾t�c���m	��ͅ
-ȡ7��Y�֡Ã]q<0���u�~��a���u-�������o[>ۮvW;cN�VƳ��Xm>38�k�r��i׸).�kq��y�ڲ�>���v1��Jp���v��'E�}�fG��{f����5�S�!~(#
�u���Ad�FQ�p㢈�wV��CyY�~RF���b �Dsv��J�[�;J���nc�%ީ��
��A9���W��{61��+E��X�~������.��&����	�LGK7s%#��g�XV�"4��o�E�N��nP[�{����Sr
ӧ��������������Ky�5]�$����^����ce?Y�Ӊo:���:��}�KwM�%)���q�n{]q��h�)��b]55�����@��SѨ#t�M�����Oх�:�����@UrN'��E�F��ٞ���s��4��ZO��1��*���^B3x!�۝��9cH1+ˈC���L ���~Ӧj~�)!񡶮���rq����\�?3Qkx�8���V�̲zh<�g�h��w�	��ea]z�}V�`�b�	�׿r%�j���f�w}���Ĺc���L2KF^xyy��+����Ki��0c����0�)ho��'����-0�H�ZAn���Tֳ�6y{t�-ʈ�\��5�Ȱǥ�_5�	��0�ȇr�2��2ە��[[�����L �Z�H��A�5"&��i#!��k'�'�p񑁤���`�������@����H7��c���v�eac�I]u�|���	1��6�18�&���*��7#u�%�B��L�������[б,0��_��bW��{�2��CBG}w2��3P���g��� �Z�MZ�U�k�L�s;���$|�(����o���r�4���w�$��́q���X���V����6���Y���&��*�G´N�B!%�rR @Z�����V��+�*F��?� q.oNÈ��%�&������i�/f��Չ���y�c�_��.-v��g�ϑ���T!��Z�y� ��$\��m9�B�O2i
b.�^�+�Te�kƠ��x�?�������>���ߦ�LP1��/��s�6�	Ӵ����ɂ�
�L�&H�k,Y�����kEO/�*C�?F��y�2�Bp�ASK������9d���lm���� $��h��vC	�B2XL� �k�u��A~���=\JJ&קS_9�)
'}yXYOK�}�7�òo��D?��(޻O�+K*OI��^u���=Y��&��.�ؗ+� �M'$B����=�����5UڪE�5�]���[���<��j� >]�S㨖4���h�IÜy}3�ڱ��5����'f/-�k��e�-�xz��+��ڪ�NaPc�:�$���M-D��'����)Ӭ8M�ɜ�t��F�G���9>�;Ug���sVP=����A'8�U�.����1	��vȲlZH�Z�d��K��� $҈��"��+p"�0]W����$��MLg:!��<ԝ:!�!����@X#��ϰ�yr[$���Q��c�0~b)^��|3�&�E(Sc+[�<�B��(�P��W�`)�,�ʡ��$���M�q��z�����n�.��-�b�k*�z.n���	2r�'�/k�wGQ��,����l��Q�(��y��<�b�J&�0̩�+�VG�/�Qy� �E��I[^{s�z�eۈ�Ļ������i�x��I�ڛ���I1ʳ��gIE�9��1�C��-x�T5G�r�.��0/9N��]aN{Wi��a�!�̪j�qn[�T,ć��2ю����ND��
O��Zr��s�^�GV�8rdo�nS��>��|k��B*	�Nl�~�ט�hf�<h?��dPr�v$p�^n*w媸� �^�v%���/e9ƒ�K����	�y�Ř�k���SE?]��	�w�d�.A�^�]�Qs�`f6���*��Ʒ�%7M�Ǜ��p�b�kM��+� (��d�B�pr*w7���`Y�za���"_H^�aF��*���O�`�p!�{�J�c+[�Ő
�-Pi�xn:�̣����W�������f���l		J	�މ+�Vӄ�vq��<Jt����m��GK��ޱZ���,�����6q���7,d�bAR�������L��RXQ���] K�kc��z/��-���2j���2�#k��8x��2d���[��mD��GEk7ܥ_�����%��Ƨ0��p�a:�Y.�s�����hzV���Z��mw[��X��Kb����n��0Y�C%?�q"ཁ@_I�z�g��2�t̗bC6Ԧ�WK?��*xM%�8찭Kڛ��q���y��(���
Ro֘�<iS�c����9r�����U���$�u�Q�5
�G2���P�~�u3/[�o�2S��fjђ�y�r�� X4����1��+���@�n�$`�@��j�����1��צL�r��LZ��0�ݼ&��
-�g��R�{)�LE��9�IS `���Ev��\�`븁'����lo3���-�s��B�"�6���i�K��HR7�"Wu&T��d����ܰð�Ɏ`]4�������L���8�+
 ����g��Ӓ̜1�C��Z�:���&�.�޲�>qP�)y��Wr�E�VKS&�s��a��7��y�� u*�SUN��K7^R�&����4�H)�7~@B��H�K4��EpK��Z���%�gB��Wh`��;�J�q��顅`�)x��w����ΚQ����v$��fgWߕb)vswf�	DmO�A��P8O�b�V2L<�p��<ɕ#��)rƓ�2��2��Jo,����ʪ#��q�dt�oi��2���% ,�`��@5�ۮiO���t����=�&;C����u��ְ3d>��i�1��b9��yc�N��\N���^���G�$��v�b��޿ߧ������R��2�c
�2�⏀4Iʸ����G�;K��w�?]���ߴ�N�\aܕ�����QtTf��O�Q����!��,k�L���7�%u��1U�����B�iK��
��D�m�@_�z>�>�fZ(c�љ�
%��Ff�߼&������7��f�a��.���ڑix������ V���~�{�U���;�\;��h�K���yn���J�MO�a��7X��qO��q�n:�yD*�6���f�1�GŀBl���Ӟ,��R���JP�Z�RTL�F�zC����R�b�*�ܩkA0Z��;2�1M�����B_+_؞�a�K�Ү]�A�1g�x-��g�����F�
�qNx�ov q�XOw_l��:՜ڲ��\�`m���p��SF�a	30�&=p��&u��%$�Ǹ��J"����LL�J�Z1,@h���'���.*�:�����x�Zٞ**x Rki@�	A��M�d��<^WG|���r�����^6J�Vw�-ӫXv�8�[f�>C�ni�����u��(�j�raEi�
�8�H��
���>�	ywt"����=�¹DIV��IH=*]�����۪�&J��۩W�%�l��sѫu�/j�t���׊%��hQ���ՙ*��z�]����dq���V@�#�r)��ts�Zf`N5c�9�B�YQ�[��:J́�x�d�"�x��B˜�mr��w#��1���sY�f���^��}��SҖ��d�u�
��z(� &0�Vf���N�m~���f�/�F,�����¼��
rҒBwb$��c�7�\rK�5����L�>j����l��G\��-K��D��G����bOT�ډ���	_�y������1��S�'�͘�*^Z趂|����3xH>�m34�����,�ޒЁ��{Q��-4�f��[
_/��w4�ϡqė�K�Yh�tO��Q��ZԒ�l$J;����pp��7UϾ�پ���ֲk���9�=9	����ja���mD���3v�b�ǥ8_��-�b�0��n(��BEq�ɾ9��,|���@�������`"�!�+��P_(��H�f\�ʖ�t|:�I�+��N��_@[���H�x�)�C���m���vg�$�T��?�ypc�F�W�����=�g0�+Go��~��PC���M��񷉓 ���T2*��E"ݷ�f��/]�:x�Y�hi�?j5?��P�:���et��ur�*����et�y�~4���]1&k
�Bف��x�Ti���4��Z�&��	��_P�"����nQ]���r˹�h�TkVH�N|���uqx��_e}�J�3ߩ�N|HCj:�?^����j^���H�2�p7wQs,���ω���^��q��1p��45:���MJ�9`!���i7h��z��գ�A^x�y��4��C�&�'�F6�[Y�Շ��b�|�n��(B"*5�b28����>����	T|Y��
��v�b�o��q��?�y�D/RgB���x�:-�=K���EgF*���Xcp�lk�sjz|7���4Bən�:ȏI�y��/[���~H)D�`��H�@��c7���V�Mhl��X�a��DW<	~j�{sxiG��da�WN�m��b[ǋ���D��['Y�Bʄ�!��OJ'N5�G�7�xY��tE�{z��KZ�|Z�G��b���#�|sǢM�?l�F�'����Z������P��>J����ᔭ7��wh���.U������ ���yo���uflS'�=\�˘nR�c��l�6�n��O�b.�<Y�$Il��֒���(���N���?�G�����y���>�6���<�Ǔ���p�
At�������C��b������>�C�">�8��"%;6E��E���f藗�q��7���)Z��Ө�L坠<q���q�n|�[����+|��
�Xa_�N�	�l��E���ι%���)r]m��1��au��\�g"��U���o�`���� ����L	L�`�_LZ�2ק:��N|�f��#|�b��O��+��E��e����td�֨,t~6�B�'
�&�?�6 �h�l!����w�=��/�)���̞���樨��_�q���㼮HA�k���t���I���Lߜu .�����[IkUO����&"X��k:2 ��@�C|�+�R�O>�f$�tM����UC��B����ͽ:������T>t��BT�H^���IF��x��%�eb�5)c������fm3n�!�N+(�?�t����]�]B�e���[�y&\PzV�f�DY9`�=������H���N-��N����f!��q��	I�큁��u��9Zj�2��Vj0>���+�~�����yq�&J��L;�d�����%�Nq��k�h%؄���b�֋�F�AN���9MTx��g^��/����Z)z��/�H%���~e]@9��߀�ݴ�����Kʣ`��	�g".�Í>G!��Ɋ��ڊ�T�}ɹ�>��::h
�pd�����qס	l����D��H�sQ���1�}2T�����eV�OX`ֹGD��ܑ����
ҟ��6�;L��=�	����aq���x�,-=����,�u���� `�p��>�ǟ	kA=�`h��8����_^m��h�1Y�K�܀Q��8�'r$�I��b����� A?wޜὉ���|;�Ȣ��������zeB��j	�DMZ�������J�:6dO9j���4bӺ���6H�FeZ��H���&mb��'6Y<_�W�C����9��r�.��0��ǢEy%����.!�
�I#6��Pw1c��-�C�B���p�zD|�eq��
�{��b�]8���G�y�4U;�Yc$KѶ�&V�x9I?2x�+żZ�sf�/e߮� ��6���;6i���`6\����Kgl�3Zo��,.N<�y9��wك�+��F�~k�3��x�.i�w�������ѩ��ܰ���B�9;1	��3kE�I=9jE�&���
��JЎ���y��EX�^�D�v�Y���b���lW���s�!ooT�����n��C�j%jY�2�K��Υ�'X�A�8�GZIE�bfW��D�΃��&ٿ�U5X��.S0��$a��bU�w�'�R��W���X����%A;��F3��ʠi5���K���&fB��G3�t��IZ���9�B�C���~B��?�;1
%�[�tg �M�c�1R@ȌY�½��zfݲi�R��\���D���J�?���B��|w�'��X^�Y1����q��ǹ#�L�X��w �yp$m�WM:���#v���"�E�ЙC?+%��1��T��S��'������N�n*���� ɾ�s����>r®s�7rm��|�B,c {L��o���l.��.�������]�'��p�2p��)7œ��O��8()��	_^ŉQ���n�"���SWhuF�*��qSN���w^��d�/��IB�2	K{�jHoJHR*��27����ԛ������O-�"��'��M>�k4$~�[�2���<���p���_C�T�uM�4r)�sAU�����t�����v�`�F�;9�Q�aV��R�s�[۟�ͳ�,Lj�c2얦t�{��g����V':Hx����ȋ��k�e�W62�c���p� (�0J��;�]֗ڲ��w�rV_IO�9~m�-����{<�>��	3O�53n���v5@_��K�	rJz�C����3���!W�ҙ�Y��D�2�KTR��4dRdQ�|�%U��CXw�`�y�KJ���w���nN�ēʡ2e�:H��� <��h�SƝ>q��;�wI��~eA��B<��mH�>�9�h�*�m��h@u��\..��>49�\k\$~X�Fr�2�B��:�9�&#[	��rK�)=Hq�썄Xe�>��߱k^5�3xc\�rw�3g�� E�i��4J��d�W0��EJT?�R��j��.%q��P׏h��ODTmc� �����.v���f�� �J�q��p�ɼ!]��ŭ��i�2)cy� e\�}���G�B������ۚ���*E�jt݇Ǫ���P�����䟇�Э�T"���a�e�1��-~�_�CnN��iH3�-���P7�FT��3�p#>���>�{r ��먑�T譋jv|+q��ܕf����v�y�5��yvg�b�+������Uo`���l�@f��1�&Mbk������B�'�l��y���}�����4Yy}�
��60]t5��>"l�9���R�H+������������|>�~_��ϰ鴬�x��#���Y!$h�sɠ�A�4�|����[@�J�&��于�R��8����$�Ҍ�>�K0��"���ߣ�AǦ���N�ݠ��3��j�h��x�����u
DV@���^�$>�hN~��2.D��v�nU�cE����%G����7�ͼ����1�|GV�H{+^����2���U���L1ɑؽ��'��T�8�X��i���gT�Cވ���ZE�m�kF4	Yj�@��?	��@ő�4RG��%>	A3d�*;^��wJ{c�^HJ��o :����]d��I����u��&
�6)P�ϕ�2~o���is"�H�/� T�sӴ��	���,?h �T�IǞwΚC�p-�)jx@��z	�8g�cCJ!��i����[�G[Ā����u��L�0��@�&;�q{�����ڝ�Z1`�YWC�m-���z�����oEYX�D��Np�O*sI����z)˒Z�`Q�#�F'J��]́ؔ��n>��@��F�%*��{a]1�!@v�9�p������p]τ�l�P�4��bK��4`7T��	��طb߲ ����q�3ԡ�V�_�<~�L�JpEh��4�5�b�1�s�2�`��s�f��c�Cg�5 l�^�#�<���9m�E}�`\v�z��T��Ȕ I奛z��u��}�}iv�z� ����ű5�#s�c�9�a�i;�E����4zݼׁD�²A�ڝu�}J������<N�ݦ��X�	Z��(c��T�/Ɯ��T^�� ���iLh��ۀ������GT|zK>T6���G�f�]d��Qq}��0fg�z
]đ�w�I�u}]T� �;7���Z'�Nm]�����%ݾ���C)� e��im<�'^{b
�z�0E:o��* ��V�_dU�����ou������Ҿ�H�Y��s�J�.j\TJ_no鲖���{�C��r��j���ad���$	f��2���^Q�wK��	t罦�'�\Qf���6��#G��R��bQOG�c��:�S�������V�+T���)�#�`�WL��,��#Ͻ�~C8H�	���>��aZ�9w��Z��!�a�����&�h��w�(x9�j���%��f����'['�#Op&��`9"�Q
���V��Q�FrFb��]6W���eh����~�
��^��*F%��������x<vi5��d��J�����͘��f����e��& ��L�v���\d�Tn�v�����C�j��Z�>�HQ�i�*|Y!�)�k�Xv�U::"z�n��Ч7�uw��T�1��Tf��z'����O�D�td�/�	,&g�'�Xi��m�|h��>�0��<V=�$gp!Nw�#��!1�h�M�_]�+V����m4��;e��v�������&@�h�L
�F��x%D�ָAHތ���r5
	��U�z�r�����0GEPEJ��G�>6{Y�b����:?�=����򴮍Q49�]7��@�xC�jrFV��~{,����F��|ײ�	,��u(l_�Ž�oǟ�����1��ɀ�q(��5/U��U��r����=b��ϗ�гJ����s�!�� �f�6������=y	RI��{9i���e�#��	Q	��5�x�l��d
I�������o��%���*�)�|!�p,�7�������/x~�]�nu=���ק�e�z��
t�g��an=�q�9�
~kU�>nj���To%��c�����2���T��ß����}$@�����	7���u�Q��BF�-�.��^�~�}��FoRy��D�I1:b7S���Oc�_��P&�e!�g�;�O0���_gj΢$������eɬ02CgYH�8�	Y��Ao�Y(�&[������ퟭÜ֟b(��lg�%T�������:	�M�o7n�#(c�_��ߗ���F�$����{}�p�*Re ߎ}�<��*���!���l |)�a1:BPs�2O�i�;)��ң�Jh[_C�����2	�;s�U�Ϝ�E=R��)py����@��&���t�Mn<��g��5��^(_����^Yc���J]�M�t@3X]\ Ⱥ@8��y�&��/x7b%z|.�IbS��������Y�2��dv�)�߭e�7̑�`�~5��$��In?N��V�а�L�UR}�J���j�/¾p��Z/J�{�)^X�D�kg	�zuSu-9zQh\�K&���_덳3D�M>�WR�u�Br�� ߶�%oo� )�$�2ᤇTp� P&���q�=2�ia�0b����)�;#����eAf�a7뿛�@���]�|p�����]��*o+(?��H�:z�����&9T[�S	���ָ8�`c�L �g�2R���t�o�����S�	ע���*m}��Lէ;�4[.�P�:�z���L���A�7yab}�He�@-��VM��W�ue��H6��_�p�A�v���C':쐩��h�A���.�*,*J�i��8�Z�Wm�)�%ظ���(͸N�����,-ƯP��E]�#���ho�Aǔ[�3��i�,} 
�BF���;�	vr*��g��^0�(�kӯ��͕0g���g�3:�G��B���~�~�"o_t�HtI("'&"��+y@"�������a8`d�zt�á��8?R�o�<�T ��x�+ҍ! G�L��em(����p�Q���,��`Lnh��_�x���G6)M��o�Z�vs���.:��K<���ʦ��<�;�:�~Jێ#+	d�Abq��2s�/>O] ��k@j_�?��G�������K�yc�ұ�o�R�Lcg{I�s�|+<��� �G��w�A+vV��
N�f��o�Ck��f(���x�޽`!O��_؋��nJ��М��5�ށ �����Ϗ����c�o'9���䊣ӿ���t~�a��4�8���O�Yi�k���Q�O��l��E�m��ld[K�W9j(��J�&MiqI�Ŝ��u2�!�����c���7�S2�5*���h&�"{D�3d̚���i�y����IZ[@,���S̼�3j���p�mz�.LF���(��!�f�T���~��{$��Vētk7��/Sdd��q@����j?{������w�������;(�rOݝ��U�=�οx��-!E[���=��L�f��zWY��W��E}�2^��A�r�I�a��/����٩3!q����֪�G!����~LEn���
d��<~k�3��G�t��2�j	]��xB�-!�kŒn��?���v�����V�똼x���|���4��T)���ƺ^����Ͼܦ�<��W{r��	�uWQ ��$�[��a�(R?�� �ɟUT�(�ḗ6�N��L�HS3�
��o1��_��K�ɸU��)�{ޟ���q��
���;n@����4���k_��Elx������&/���	��.�⏛��|��q�D9��!�*�g���~b+9��D��r[uW�73�ab�F5�$[7�� b�����=0u\ZB+ҍ~�B��cK�ۈ��˸'�k_�h>�W�v"zn��D.l��]���H�;Ef�k`r'U�mSV��q4T]x1���G�}���桥U�L��;c%2��`ւ5<|Z�̜ڇ�$��.@5� I���A�����+�$E<������j�=��2��8�#x�x=(��f�R�n%���=��R�(��[o*SU����K����eQǿ�gA3ON����`O�n�uQ��[	Qy�M�9XC*}i������8��S/H�dFYr�t*ၻ�t~|K�n�J巵83��x��ꪼ?�#�hk����s�� �"��0E��τ����1�nqs�X�\�x�oj=�e�x6��p��������V���s8Z�:Dg�'���K]����}�W25kSR�=�Nb�����u�B�AQey���?�~�� ?��ϔ�~,;m��Ћ����Ԋէ��n�! >�Q�)��	�G{SJ�J_�4�X\��+���YMap̨���X����+W.H����tp[SY6��>6�>���rQ��w�&�J.��P��-ڞ�x*�q�Q��M+�Z?��
�Jf�C8�T�v�Sn �AnS�}х����;�\�(�oR�+A�5k�����\���E$ױ�n��Mx�6���F����$iOX�L�S�6��w�n}��t�F�sɞ��XVg��O0Vg419{���%,��{��B�xd�gr��A*��@RF���a]֝r��HwIh�X����γ��|犯V�(Φw�/�(��g�J�`���Y}�Pqh�x�jb@�!%"`���Xs�$~�]QHhkd�.�	$��R�8�ܝQ��;Ǧo{�+z�NG���My�uK��V�oz�����%u8�=\4�د�����
�cD�Z<�s_hg�}F�p2�/6GO!�9�ʴ_�[\DA>�2����U�+��Z ��V�`=ϻ�]�U�:�ix>:c���;�l!}�}��.Lq�/ޑ�*4|o�����"CC���TI���/�zV�}�I��9�
�8w���'�.q!�'r�]>qs��R��S�V�R� �BC��G�l
�T�H�/B�Z�z H_J8�+�i9��D:��}�u�6���$^21�����J_Q)DE�c�_�3whݒ���O��jX�A<f �St�S+q�0�w�O���n���h��@ץPb�l����4�8���� Zu�}$��H$S
��2���U\��[8q{#�{:�C�W!rAC�Ӗ���Փ��o�.�@��l�2��ܱwfT�J�`#zA�QtU)����2�"'H���Sy$�6;3���po��_~=���*,��A�l/9 ћ�A������W�Т���G4�D�5]����fw��_hZC-�蝃L�W���W����5��M����������M���@ٔ~w���D@��S� ��� �pω{�r���\f�xW���-A����N��vqG�|?����b�7��-��+㨁u����.N�P�b���]~�0������ö�G����o��!U�[���y�>p%���dТWM�)����3�vϒ�o6�z������j�	�ODUS�Yt-�y.��V�w�I��#�YP�%趙ٹ���O���8����\Q�o��/5@S�!��Q���p�Aaw�ތi_�g����N��ȥJw>��c���텟:�^��<c����}4�[-�s�wG.P(�H���Z��*��:�����3mCo0�eh&�,�����Q�l@�����l{h��2�&Ҵ�s�6Ao���(ϲ)����wj��)�Z���ԁ=�'���������C��zr��2@AJ5O� wA�&�\&��QD�&�{so	�fS��1���h��@m!��%��8�"�W�Ձ�H'��t��5y�3(�}w N�$i����7!���q�p�l��Kd�������y@chh�
�~g`��_��T(�r�V�1kz���<�k5v`�X+����hHL�N��W��O��.C�l���5ZiD/����v%23��Y�"�?W=��$��;�G���nL-� ���
��8U��/ {)@����_�m0���%�MaM.��Q�l�Hھ��
�haSA#��Q�S�N��"Eh�T�y�f6�Ibܥ�_�s���c',noE��g��;t�K��&�RѴ���x�E��+��k@%������-U�ɃڦG�W�u-���P�כ,��
�Ҩ��\�m�9,��!��zݼ6@M_��,�V��e��+s�	)��йTdyd���
�F����9����m�"J�����
k�ɜ}���RUr��5{���j��k���	��Ϩ�~aB�?�gw�:��؝!���5u�z��a'��1r:\�C�*�e�x4�{%��%^E�����dnA��y�fb�@�T���r\��}s��?�����M%3%E�'��C�*u2�3}��k�o�s�>+�7��� �,����=!�`�\Ad��߁>�ױ9�Q�E�D\�1��v�?C�HPMĔ�G�,N!�`��_1�������Sx�Pl:�c�o������5^+쑖� ������T�2)=ʎ�	t6W)��`��Y`"�s��G��^��T�:2�cb�Eo��$2s���-��$�u③�B�Nz�W���(%1#Z�3<���n~bb�8�r�.I�F�T��Hz��Y-tF�EY\0�]�g�Xe�l�������h��,P$n<���ޏw/��o�}4;��L�f�	��M�%e X�T7'�QK�!pL�b{��s�s�Nf��Ôu߁l�ʎ>�U���@���z����H�����b�<��C����]|'!��}��+nR\��'�bi�4$|�v��J8A���}����*�UrvSsi�����:k���BE�6\yI�!W�ߦ@�;۾������+�Y��ӆt粎����Ǎ�v=KGs�#��؁��kJ��>��X�a;?�������L_n�3r"���p'����Jeu��ţ8g��M�p@BT+��}��L:+�7��]�P��v:_F�����r�e�DIT���C��D@�,xh�i�TJ<h<Ǣ�V'J�. Q>U�qY��xu�FxA�̔n�*pd�u�W]'Ƭ׳���È��@���{a�����xp�Jo͎!]��~�3i�>�SCĥ����c +��A]?��V�--�9���[s�c������lFh`�]m���n�}���Dƫ� X��q��mZ�9B��U$���6��~��!�y>j晏|��F�\����Y��HI>e��:�_�DG�
j��M�%Aʎ��������Ǩ0(P��@ЊL�5h�%�(r�%¬�����ل�ȣ�X �۶�K�U����=�!�y��M)���X��@�z�U�k��B������L�G;�P	�3)���SH�����*F���؜�ò�o�ql���^&+��
B�7���jT���M=逫%gUg��0*���.ߨ�K�v�F��-3�ʯ���ELuo���r�I%*�I���Wݟ��{l#�އ%R@���щ[�I�C�J�U�u�3�ؙc��b�d�������#U���=�@�b|uojP�뵞��2���#�\��͂zmK+8�J}��	�X?�m~>�kwF�#0x��;]qWUU:��d�aQ�����	&5V�?��v$���<�r�����̬��b��x^"¯L8��������Wش��C���_�MmV������6�/r�J�U���Gzy؉���j�ZU�yb���qG?߃+� ��s|�-��btJ�޼jE�`���û�U���-�j�K��TV�W	R;c�Ӊ��聩�ǵ�D��~���#"��7��Nө���q��XP\�Q�
�O��V�vI'~��6A��V�����fa��h]��@���u�U��iAC��p[�9�l9y����K�J�ƥ��(m�Aj�rA+dX�p��JT�Y`����"�\���h�7Ee���.�-��?�[˰�1i[�j����s_�+�ON�7>L�7,��T`�?tk�2�O�d������.c��8��c��`��<^G����љlX`E���#q�T%���;��Ӆm/�`V@�~��<�=��sN�ϴ�O��r"e� κXIH�,	��u@��霙�Z��Was/�2@X;�Z��Ĉ;��4��I0������:U�0�W����U�-5]��o֔Oգ��BR���]σkd�b�}���烦 #nmZ�L��l�A�0�9���C�Qj#O=p�,2���U
�Q�Z!$Q:	827(��W��~�X,�,�"L�ܙ\����n6�+<�	
�=��,�e������y�����¯��w��������S�tk13�2�N5��ԩX��u'�n�1��}�ַ�~Fw��t	�5'42 'Z�"DV�&e*B��-@������,�e��9�Ѕu������g	�q#0���q!#��f)Wt��I����9EҐ\����
�X�R���jh�I�2ё/�	}�(�;
B� �7�K�P�τ�f��iG��}{�D�'Q�Q��bD��rz�ϒlm��k����h!mM3aІ,���h��<X����h?�c������o�]ԟ�d��e�M\mk*f���M�'
�2�;�+d�U�,� W�Om�hR�M��Z�k ��ip����C~-W��CX�f�Y">����|L=��}�[O��GT�q{l@�Y�RGW�7_�c^���D`r_�8�rV9�)мdn����9���l��[�.ln\#�@KN��"mr����n��u�)��Աu׮��9�*:7�(��{ّ�W�B1x��	����w�}Q������S�a��8�t����j+��\���������-��2oN�2q�? ��ۜ鋪�����R�f��wI��vN ���Y�k�γSM�,�#����M�*L�B�"F�[�3��;z-,a�TAx��1L��9r�0 ��Td�B��_�K�:=�	r�Z5��`�j]�w!���x�!��R��ȽV'?m��m��<��c��Ʊ��o��!O��/b��'x��w@���1��2y����ѹN���3 �Tt��(�0?��Є�h3�X�u��c�N�	E�Ξ�=��d	���ώ_��m�|y�DŬ������EÄ̿C>�����X�x���H��AQ�`X����{���Pu&��PE�u'!U��\�)��묣֝��*��?i�u�@Fȩ��Y>�����(䭅ES���<�jzҭ�IS4a(�ߒ�a@K6+z/���4;�e����pe��wU��H9+wk.Jl;rm�L��W%���p��q�{���9F�@��8�\q�+�E�n�۱H����N���D�+"��g��
oO ��d������y=[v�`�:2)��T1��y��/N�G� %ҳ:�b_� �Bh�sy%<�%wl;b��ԡE�N�u��ָ�P�D2C��A*\{�!j��6�Rl*��;���������־��/�QƱc���:�L�\�����Vu=�zm�|fHӊ���ᤆo�V�;�U�ƚ�`�}m��7c�[�F�� �'+ܯ�o���iwSϽ�ݑ�r�篡[�������F�^�QO��,����:)�+�����;�B�@��#Q�7��G7"�ɕ_��w�����2��'�v�-��{�j6��W�T�ng��6����J�P�^Y6Z��Dq���B��j;�����V^��i�ye0vRKr#*�W��MFQ5�*$�rumA�
�W�<X-�<����P=$�����R��$T���_{w,�	q�y0@n7P�a���yD��y#}9@j�v�ösWߏ���}��'�)����4�ӻS�U]�?���<�l�p����)1�QH�"������c����ܫ��i����ǅ��(9�nS(7�|��6�X�w؃Q��7s��`c 쩃8�Jizt�\��
bN b�Y.�?DxQ\��4�U.۾����j����p��XX*Qx�5_"Oګp����n�a�B��A��H?7���w01�Z��F �-�Ѭg�FrǢ-��
-���#Y����9t���V2�8�Ho*W�T����W7������n��l�]�������S�g�}"Pu�<GQ+@��$������zU�h�b�x[���N)���/������s�����΄?����\��~�������L^V�� x��w�.	l��hQ�irq5+ӢLC�c���o�d�$l��'	�Eի%D!"�COI.v�h>4 �.�i-�v�\��V��v�O%�$��"�4/]J#p�_"���<�{Y�����ϢFx^�rR������	K��>��X�G vN8p��q:��uN�T��p|{;QH�D�PR����*M|��a�v��15R�>�h��E�Q<�PP��<Zt���Hl� ���ӑ
/��Ѯ�.��=d�W#��@#"��݋�/Z!�L�<�[5�x���]E:�[�:[��W���E��}�� V�h��φ�/����&GK#�!����������sU◥-,�'�RZ\+DT�Vc¹.t5�{.��'	}j#}��~ď2ԋ�������5~���k%ap��F��q_%��R�u��NM�W���3�(�����e�Ӷ�T��#��4y�$����T}ıRe�(`��#�P3;����j����V�0��n�g���&�Iv�~�V�Y_�
QB)��檕����X��,�L0��.O�l�i�aR-��O�9語�) Keq!���7ج=��� s֩Am٣&�ڈ�0&A�vT��t�KDi+��S���#��T(��<�ń��~���K���̂sF�m��Q��p'v�Ü_Un�����ecw��Ԋ�Eэ`:"J�L�dҶ�9��y�2��~��lo�N*0@�)M'���.��5 ֵ
�K$��mPhR���._5^�ͷW\�sm�j�Xu���Ub�da$\w�$)���Q�W�����\ރ �5U���1��C>�-�H��]��u���dCl�]vSS��)b_��3���J��O�I���<8nb��x)�Vx�r�@�F�TTx�.Ț2AH;�·��HA笊�Q���PPdGm�����b��\�Le0_'��#C��jg_06+�I?C�ϔ��Q����s�(���f���'Nvk�7�9��@�{
 -�|8!ȭ������,����n���~V�W��eX ��~���7C���s,��Ƙnލ5�Q���=��&�&�\����h[�����L�?��p;���)�+��dg�ƨ�������;pU�n�rn�RJd#�E'�ZIM�c�՞![��X�V�x���Vz�#���8ޞ��������}&֢��"���[=��@ش��z-T����V��g��p4>Z��\�J9&[�#N�R����1n��1F���PL.��Jx��o��JSz�N��×��V��Ձ�[��D^�ν��r���h��uhO!��W��M�?ų;��o٥A�z\ͣd�@U����v��>1A����irV�b>_�fp#�����}d�Y(����2��� ��{P�밸C0_f>W�d�����X�h���e��`���(QQ�n�ԟ>���;qT�N�mdG~�{w~�!QYq{߸[O�Y8o����;+�����=֒��㚴9;���D�j�������\�FW�}��P/�@e�?4���_§n��h��l�a�׌VV��)<��W����*.��Rb"�t���P+���u�8�+O�J�5���s� �`�_����-I M2��5b�q�_5�4�b�7p�0����������"�1����%`���?k�M�Ӈ(�WU�mQqP'�,�r4�Β�e��c6����W�D�Mq��q�z�QP�, �E<��T˒a�X���81�;~ )3���_�	���ױ_m���w�l�P�H.�]~�Ȣ"���������� L�ނT��g2g�����=�њ�`�ظ�m�d��1��o~�9�~s��F@�d�)s�ŲX�v�<-���uJ�K�������k�)���<�\Ħ���<0_�o�$��v��m��d�����r9�t����»�L���x�GɄ��	޸��W�eϔ���(��b���'���ID�L��y�,�ܞ˥ňc��l{���%�@.��tQw?�Ĝ�Q�+�Q믩?Y��)�c���_�.}*�zTfB����a
9��n�s�{I�-)�aqw����ݹwl��]\��pт���6���@�H�Ɣ������.�^�ho�,X����z I��L܎D[(�Xb�Q�{�A�_���-�� ��_\�wW��
4:��E�J�OUmD~y�M-��
�7����s���?�����D�Q2�3�Ek�y�U[�W!��1SoϞ}4j�e���Ip���}5 j1�܉2�t\q?�����Z�`��� /� }�O1/�?�^E�a8yA#�.]���qz�)yK�S�i-�o��������_��It���si�*
�nz�1Ձ0w�:�zp�}Q� �����^�Ha�֎"�*�п���T!��U��pOh=� �� -�A�zODb�"sEԆ.���'n��*4�nȑ��q��$���Gt.�X�w������Ǩa�=R��)�{[�r2>k^&[��AY�ą��4�=\�8[$��WX�R`��SJ{�wY��˿�&q��� >W�/k�ڱ�nc�_�7�Qk2���֨���ʫ��BR�,���KJ��E�����l/cYש�n;l����}���E�F�!ga)�OPe�C��{�^uR)�UsRX���7�w����7,4#뉅�����)�� ���	,�P~�̽sEaE��w��T�V�����!u�I�y�s����	�,�~g*���[�MT�p^D�����e����@Y&=o���Qk z����ܹ{����Z�
�ꡟ�A��]�M�q�!�rʓ9�$�XCW(��?4h�u\������C	^_p�Ն��@�ˇs=W��yY7�@���`Edd���J�É��4F���p�kr�w�_���s�o@E�l瀦�Zw�-���i�d|g�M�c?��%P���9u�Ή�,���_�e~�Te)
�2~L?Q�����g�P�B�waɻ'Ԁl
10�ڱ=��-�
�U��d�cDT�?ރ
sFD��Dg��z�!�P�ܜ+��D�l����8)���׎X2:������/��]y�ܘ��˛���H�rRY1���B"`�C�͎�'d��#脆��P�~�����p�?qH�Ns�а��j6}��ڗ��+�J�T��f��eޢ�O:�w�b(>�%>ϐ8��5�|k� ���NkXV�Jo�C=�q�Vwe
I�=3d�?���Y�����JG[(��<�O~�w�ӊ ^=��@�y��l�-�3� C��9���m8��3��/:�����x���s��L�8��Ef�����`/��UCfc̘~Z�/�O���a�	+.Z� �s�Nx�N��fW�=^��W�F�Gk~�(F���ݚrC���v���ӝ�p-.�M��܃:Vt�:�XP�-nX�����<�([�9���� R΢�}��t�˨�W|0������mhC�{#����b�I��e���tTs�L�[(����[�T��'� jr+%�Κ��N_��4������ւ�e�K�B��J��b�6n�|��J�d��;Fuл_�Yb�Hm����ޑns�N����P�`�BĴ�?�r�O�����8vE����^�{��;W�H&7V���)����Y��z)S��p��@�zN�gr�d�0������j�ٛU�g�)��Ӫ.9�!��X'u��N�����rUc��Bx�oڻtN�Y�0�������_�&jʭ�W ����"F
5�iy�ٯ�(ԏ�:C-`OѭJ|�t��YF�����/�W��g��{`yw�1��,\H,m�f�A�}�Z�Y� �z�C�C��s��Ir���q]u�R����R-��zܱb���-��"+IgPފ` �I��]MϾEw-���U6F��&7
����UΣ�0:��ў����֮����qq �<���<DM*��m�����H@�w蹲��>~]+���P�e��cvz/t�!I%�4R�8�=!�������Ւ�q?�Y��n�kGo������ך��gm�Ʌ���}�mx�d��λ�z^�}��F��!�D��I��B]ޫ�Bj>��w���P���M�0�h�`�'�8�O�����z���ׁl1O0C�(���Ҥ�E�A>��x�`��4&��� �E;���~�/�x��J;~��j���ј��0��>'��+]���'$��c�a�b�M�A���ie�-7p��X�Wb��fj˪�+[�cH��%gMir^0Ar:�x��I1�� �O8���0��g��}9?�%�7@�  a��SP�H�m��q�$,WT9�4Pl�����5��!�t��ˏ�:����H*���`GI.�X]�{��u�E��c�����{����	4�cw����q��9.vKf��t%Y
�rZ.��b��"���>j8S@�ZΌ���w0�mzz`�mr�+���pSy,��v��Z��<T��x��-gd�h,���U�$i�^ۮ�R[�_$q�y�͓p�)�y�c�#��Lk%o�gg�|�m2�?��20b���s��F��{�E�a%��ձ�(��Pk��I�tV���|��	����A9����ٖ{�P���jC�I� @��8�6�D&�O�V�4�kֻ�8.α�
	m��$����쮴��+�w���8�G-����ǻ�Q���}�z̏��k�E���*���G� �s��r�Xc�D���S��%�+�C�r6�wP�&+�IJΈVfz�[bC#����A3aqJ!�Jzg����St�Bhc��>ȑzj#f��'J+.�:P�	m"^W�	�+^�e�'��ay�k�ݓ�O�Z�"y�׸ը��^�`��9��w՝c��dt_���ک����e���l�˞�����z���tv��S�XO�b3j��eW��BZ�BO"����<;)c��# �\<+���0���pHbup��u_�L����W�w����Z
[e���
�	�~���l��=��w�u�5�I�Le���#f9i <��Y2E��K�_oz�)�|&�~7�?k���v�����
��k�:�3�sa?RKR9��rTm����~�t;�q�>��D狒x�=?w�i&�ՅJ+�0Qp���;ӎx��������A�ѡf�&F��B�0&��f�x�K�L22���.�W��Ʈ���7'lg�2oP��%���TTK0f�!p�ݏ	��c�l�4�e�%#P�۱�I�)��r�R3���� ��X�)�Ҡ���CVև��jv�˼��ޠ�	CJZ6֛qm.�;���7!D���CN<�%�-�=x�>�nG�>��_]ޥ�<�Au{j�m����v�MW�J���e�˂��(���� �'��	n�Т��%�O
�p:��(�${�� ��P�?�$T�?��_?�,��t�4��F�EoZ�n��SƜ����3�6�U�2vO���Ŵٿ�#��Nف8��ƝQ����H�9�U�&�z3��ǎR�s�=���9$ё8����_]�F߾����U�2�{򅊺5l����9�7���7�A�ސ6����O���Do�
�25`�ܷ$yJ��蘆)�e <���90�R��wd.��e��rru�-��!0�O���A���'d"��p��>.�_�LSBRh������e����WFX��i#��>�a9wة~3��N�>��x�Z_0"��}xN$�o�&�&Ec-ߎ��h����8�nf��:b�J�!p��	�s?�),�¯!RK�aҦ�3_�Bl����_�63���Lht�N�ުJ�pQɋ��B��s�4p��P_oXuY��B��!��3D�Ut�A�-��>l�H�����nW�oMU�[���[�Rv�F�u <��q��C�-�w�=	KbS�>[���6�M���@k�/q�oqA��m�ڂn�ꔍ���9�����նK8��A��0�#��u7��<:?H��h�C_�0����=L����7��6�Y5_��Z���:#�C��s���ȳy ִ遦kj�-��>9�}�qVe��D�䌄~�p���}OH�Y����C�󶟤���{�
�f��^cp�{�G�f�#m#d?"�<�����O��	�蠔5�U����~�U�m3{�]i�g�,�W�_c��8T���	��.�O�1�JM���X��c��;�qz���s�]YA����˜ƃ	qp���Н��
���sDS_^�I�:|	T�X.�lʎ��J���%�Z���I]����C��a�UX�Թ�G Uȸ�y���S|�ل�Ud8�؄�Q%��Ni�z�bi
%�l�өnS�Js=H(�����ٲ��~U�dSS)�T���n�YXK�Bs:̂��Bj�~����;`r����R=�B)b��9BE� �hj�B�@��dN� ��CZ��jؓɵ�&��X���D�L�@�d!{Y�ş�P%s8��51���o�E�d�����}5as@#�Z\�,�V*�8*
gO	��0)Ք2��35ɳj��`zzG?�ֈ�؈~�=��=��i�ǩŧ0Ã���=�no�胍@];�	�Z7�c07���T�̶(��ݝ��ɱ'�Wm����rg�A� �&������*����+��%&����:�A%�q�xF�]��81����lF�qy0nr�u�@�������+=�=����~v�|���D|�d�62�+��t�֠E�q_� ��Բ U��tFp���W*q;����#�Z�N�G�o�V�UT�v՞vy9](i��V�J�J�_����'P�w����Y��i���;��n�:�k\f�S��s'n(a���)����#�2��r��09�]*�;Ӭ:G*�=�s9Ћً�x��Bv���AX��y����3|�uw3������3����g��%�B~n�Dp< ��̛����]B'ⶎ�F�!{�F�-C@�ښ:�l��-Ny�X����j�?��:���{\W*�^Q5�k�S�'W}���~��}��ኹ��}�z��G�h�}I`�|�پ�k(c��]�K\*[4�i
�ق�@K4q�����?ZY��K�}�~�1�4���Gn�yZs-^+�g��Nd�#��H��6��;=0<�3������F�| Kq�I�v��T�zv��~pζWW�w��T���"W�:��U�1�C���w�?J:��ʆd�#���*y�词j._��<�!���3r����tԱ�.��;��*����M�To����P7�}mŚ��!�����%+"��o+�����;R��7P��Ҙ�a����0�������g"t��Y�}�!Tv>aIB���/� EZJ�  Ԋ���4J����w�3f�#�S��Q�`� 
_#w�����NT�)`	�=�s�m�� ic.`K�d,V�~'�Ԗ�d$�N�����
W����fIKB�s�UӡFʽ����]#m<�5�[I��#�ذ��k6����3�����>܈�DO;�<�6x��x�,�����a���[y2�g����?��aŜ��Wz��|��1���xUʾ��/��h[.������H��e��)���g�#�Ӟh�#�7��i�[��.#1�c8
E���W8%=�R�	��2fp��}���d|�)�ݍ t�.J�&�v�z�E�8e�u��?7�ϐ��ws����~�}2-z�Z�+�qz�@�O�gz2��L�R�ߖ���i:����`�i�j.X���m��^wDԗ� � ��p�7g-׸��A�ڃ�^��K��k}�q뉼�*)��i�mh�X;C�b~�9�/d��9kZ��0ΉS���>�S}��01�>���}QIX*����lm�L?p]Z���,�w] ��w���CF�-�91�ͻ�hu�I� �N\�GjD/�z~����>�A$\c$"^^�K��6yO��CK/p�#li� �$�`΍B�{����I"��NXTT��� h��5�%/g��kwe����D��Y�h��b ��l���:�(�ú6�*H�w.-"�r�rd؎�cyo(L�\��̐�b����7T`��ψ6'��)�`�������HÂ�����ĥꭤ��*���`�R�[�ŉ0Uv����82���@o�ޜ�n�0K�"7��҃g:cM:�suZe�a
Mު�")OF:-w��l���o��v���{w��+B�RDTǛ�-��c4��y_�<'}
��=��!����Џ?`���
�洉�� �V��w�Κ9�˘������iҹ����A�
� ܖ}��N�n��(%Oųga��Nd�d�ſ���_�4P��.��v=Z�º�����:;e2<w�
G�!`O��V��6�F�
(��	�A�T1�
)�Xº��Iԗ�vd������u]�@��6W�F�4����H.
ZA��.j�4����)TC�5+���K�5!0-ͯ��5~���r�M�[�m���q�~LA%����2~�yky�=.���8�*'I�rk�cN��i���}=#&a�`5)��qb1{p�*��i����8���S��r<˛���s�����>�������g����?�Fʓ;�JqĶ�M� }kf�{�\1���S�Ҕ�BJu��.Q�kR���O�7�VJ���^t��b��\�@v�{ɯ��r�~"���!�
nx
�
.�?�U�������p���s�{���z�J�5��p�VȾ�.�4�4	ચh�Lkp�t5@�hDpHƕj�ۄ6���h�T�7#j^�9��X����i���YLҡB�m?	��<:k8��°��<�������������FK�����O��7��VË.=r�~�J���ߨq�l|p��%��u�ֆ��N���9�w�hs�o��Ԥ����>{X5��qLۓ��S3�H�=��TÍ����e��6O����Ǝ2����T(��6�@X��B���:��f&Լ�Є\B�l�lEPԕ\@l�{�'����$�?iʹ�߉2kV���(7c{{p�����=��m��d�e��Lǌ��GIGY6�\��Aw�%�T.O��ľ�K���ݪ��O��8a������*��b�?�*�tD2��[i�Yw��m�s��b�g���o��-:�>���'G�9��"�ɰ��������wh8�G04զ������ؙ1[��Fg_�Ť�l��)�Hc,!�U�XP�L���?��-�L͘���|��C7#�Dv����)Q
RW�Â����f��Щ͞�h]|�v"��MDĦD߫N�א�h���Z&D�?nc��mѢ׍d5�h�mF7��5�L��y�b �xϐgdI�.4�v����u���]3��O�gK˲��"]������@PW�i�xͶ�.X��gH�ot�͡�\i�������A��P��M��c�L��jI|}
�2M͇iA���!v�P`���h�{�]���{k��N�����Hͣ$�]��.�e�Ǩp}�3WsO�6`���	��چ�f�̧ES^�^s�W�����-0b@r����ʾJ'qG=\,Z�n��kRl����?n@��a��B(r�D���k�������6cc��K9�#�n�P�E�H*��W +�����,].�[l��]`ro�3r�뙌.��I|�k
/���x\^y5���s���v�K�<���l�:�o�c���g���z᜽�D��4�~=��rc=&�o��l!r�����f�&:&D"���;I��U��5��{�]}-^���x<C6h̯�(Ħ�8`s.d�6y|)�S gBQҷ3�ew�1�a?a�A/�@}�����O�/[���Hl��ѿ�>�����Z$�'��Z��>c���w�{Z�&�):־-��\�Pċ�r��gڼǋ<uRW	#v��H.��[c�r�1���S��)Zπ�t�H�� �~i\�w\� �w�c�(��P@Wg�.X2��#A�`k�
���犓.�V-�O`�Ҡ�7���'Ͻ�k�q< &�`�P�1�=__L:��qR9���[��������)
^�͙%���{!�Ḑq�|T���p�5<,=g.���?���Ԙ��;P�q[�j�2Sk��twF�1�G䨅X7R��3r�7 Uo�g}�8o4x5#��
H�w��#RkpI;-����Łh�I\(��O^)�NMysXV1Ԟa���Cc1�ڼ�qA1�-9���k��h���SQ�hϊ{�t(�)��,Na����lt�B=��)Y�2Y;���]Z�/,�
��V����?�7*���X\.��O]SC�l�)�}_56�"G� Xل��� �dų��eS�����QS��������o>n��P� ��k�q�Px�x-ס�Q�8��A�̻tF�qqaU_����P���(H9|'z��g?��Z��>��ȍ-�I��t��{²�+i[��E��j�B��cZ��4�״~/��y
0Qw�s��]���قQ�Yc�'� J}=o����wbw��}�4��S��ҭ��T�!N����my[����ݩxӒ�)0X_K�BSʗ�(�����wQ/5��N��>����77լ�s����V���_�(�D��hp&�Z���;����R�^/{��3�]����{o�a`|�|��+�8h�)+%Xt���كZ��G�]�9�8h##*�8�H�p�O�H��0H��>�ry�I��!"��U�?�.%TS$����菕�δ�P�?w[Rf&�;�����yJ�s�K���x�A����P�=E}x�F�A�
����ؓw^��Ӆ0���:�}Ӆ��N�ڂ@g@N��f���%����}���Z"����,�6�a��LL%>K��W[j�u��������E�]U���?��{�q��u{�?��c�D.��\,3(O����嘅�����ׯ��1�E};�Y͑#ey5w�,ڮeùQeDA�D����A+N���q64u{����O۔-Ѣ�KpV4m7�~d=��������Hw�6%g�ς������ u��r��,ι�N�NJ6�jm]��}B�[)�nH��p|X�Lt>���^�m���r��/vZ���{�\-IШ��̢WS�X�e%H�<'Yn�fRL�.ԥ������&���6��`z�{1m~�iI5VA�s���X�S���:z Bu����	'�T��mC����"���Hj�KN�<K�E�gzػy��ȡ�ڋ��mAwk��ȁ��ݱ���2;�ʹ@�f�i�fM���~�����^�e!$~��9���������leG����2� �w�Gg���tT��?L͸:�Ri�����`�.�L�e�u����
��	a�-�yi@�e�]���l���)��D���0d[�ϩ*�~���sJ��/yN:�^^kaAng:�9�lQ}7��y�R���8�~�@�l�xC�k�)���!}������qJ(S�ص}��l���t�x���i�7��_W�����~_��ｈ�*���8d�S�0\�A� HYx7:G\d"�Pϟ��Z�L�b98�]�P����Qk���蘭ԃ�:{��'��޶嫌N-F�D)P#B�BF+���ݒAxC����a��{�T�
�Zt)y,Qz�f��|��L�R�Y��_���z��Ï�.=6�WЦ�?�㭑���R�{p��7'�]g�d��y)���x��8�Oo�ni<J{���?���������U�~}F���o�� M�4�rv7'��`��B�������"�	��Q/����e᪐۷n'_��k�@�0p�~!��,H��/"��X8�aD�b��� �]T��Za��+�$#�H]��9�}�ZG��ҷo�0z��=}����g��W�z�洍<�$9�7\��𓭜՚�c$A�Ѯ�8&�zox�@�����H�ȕ�c��w�t�׀rv}�B��СT�Vt|�y��4�E����PWE���%��s��Uܕ=޵o Ħ�{��˧�!Y�G��v͒ص��Tw�������Kw:ċY��+&����}�c�,=`5���E��w9�)B�-Z�m�"���#$�=)K�#M:��	hB��)3�L��˰�vI4.N+�</���=� ?��"��$sT1+zR���y&i����+�L�Ӝ�d��[���+c`oh��OU�nK�8����y(�awII�ڏ��?�F��;i����(�B4*�u�QN��B�3U7��"��F��O�ȸZg�G�G6'����!{�H�Fs���V?\�W���w�T��u��~�1����:��7Z�\}Mr��3HT�qXgS"��*�w�=͒�E�o����7��i�n�h*W5���\��R��o��#�AO���b�my���_6>�i�I`�!w
��IP�5.i����P�C�4���ò���_����ϝ���x�g���>��F0b����"`�_ACj<�D9�t�r��,�3ւa���ӥr���_Ipp�����i���a�N+i�*� }^ Ω �Я���E�|�>O��@���k�Rfێ	� )��gB�
Қ"V��h��"��ۃ$O��۲�W�k�wO�ԭN${&�:�)��rf7��Ea��P{E��k���bV��"�0R�*�ǠE������	�n�f�W�S }�4�.�]�D�-����D��.����#^XGd]ChG�����������!l!���V�h�z��&g� V�R�HX�~{W�N)u�[��n��k�t@'h�Գ_��o_�]�j�"H�2���x3`����>Y�I_zZ���[#e.npN�e"�h�<���)\�f�+Wф��g���[oBҀ?P�s�����|?��Am콾X�Lm��{6̕�9�A1aZd5�d˯���hס*q�K)PPH^AC(7� �����?8��|�y����H2�����=�60
'薶�_l�Ur�ri��VS�K4c��J�0y�&�u�o�I��m7^uY(��!��jB������ۉ�.6���R�-����� ��	k�ߘ�ć5��(���F�7�A����>W��i�TD@f��~s��I�C-��]w��zߺ�W	�g������m�/
��t��
�c9�)�͉@�ԛ]�)Wt��׊��F���u��Z�p؎�0	j�G�0��o,���#r��@�ˤ���+b�
�9��_�b�=$q��k�qÊ�Y?�t�6S�|b�����_�j���^�կ<W���դ�8sB<��a��C^��=ݤ&A1Y�=�tu�r���h&E1+=<�;o63�ƶ�_��ڥQ^������!Cdo6zї��`�^̐RTmD�L�2%�sG�`���ʟG�_�N�Ψ��ϴU�q�X�_�滒�Z�����tCgN�U�te��t�;�>�X�ڥ��8������kZ�Hj�Ȋ�ͧ���|���WM�B��Kʗ2=���]􌍋*���~����2�>&XS�Mt��>�xX ��]m�����o�E���1Z��s;�D�zʓ?`C�*H�c����x������D����W�D�`�Z|si<��8��cX�3�����F���S�>ػ�e`F�'��|��	osѽ�x���� $M������5>�V����C�eB�nK2�� ��n-t�@�LX�4�VD�Z�t�m�T�m�mz�WHW�_;o�=2����� ��U9?(В�+�u����U]V��IB'�R�Y{#��L-*5vH�A�D�`���Š�3WZ�~�.��4.H)̩�kI�n[��K�dUƐ�<�%4 �H�E�2��ZC�]_[�-�Ld��8c�&P�͆I&�>7�%������tq����>nj�)Lۄ��B����R
��>�d;�(�\��_̭���"Su/K�K0��;�m�������h%�����d��Yg���E1ꌰ�s���3-��f�)�o�3�T߳*�% E4K������lݫ�_i\�6��tޭ3�t�^KD�9R�~댚���L�� �m�����ըo�Eg���~'�+uj;�����2�^�X�h�'��4���1Y16,cݶL_�*�%i
�^����u��K�@M����}U�w5n���1���Ȏ����֌$��C�20�#�h�3N&��4W1Z��� ��L���a��Z�P��墙w����k&���u�XT#�T��� @2�_˽�\�(	���W}��Ǔ��rLO�J�����������l�l�k��p�u������A���$��؁`r4���j��H�!����o�fe���U�*C
AS����=�V�$1n~���a�_�i��dK�M�r��/'���ArB�����a�4Qr_���W ����i���\+�Mч4�Y%Z�m�H�0�����9@r�mL��dqv߲Q�.�jmv�^E�"%��r |�>m��~�n-�ULB���J�f�~��������h� ���:�t�&<����m�ٍ��]��ת�H�Nwb�����Pn� 7k9����̩�TK��B�f�d�S����S^Zx��ݭFuvD��a'硾���AN��?��?�V��<κ�i>�&*e֏�Ē�0dJ�s!m�eB����b^/l�����Ȉm
�Pi�3�����4�+
��l����=֭�3+VQߢ.��:�0>Hk/w���겟 ԣ�*N����S�ݶA"ؙ�������E��l[-�LL&ebɇ"7˰���?�}��j��Cn�Ɏ;���/fh�Jo�0<���<ǈG]K�T��k��%�1۾ �!����>UG"a��m}Mp���R���]B,��Oݤ��:����3��C�	�{�µ��ښh_�u?����P˄��:�_��o��o�Z`��X<�$<�Ҙ�r�,p�d;����3ؘx4���99a�LV
NFF<]�����Hp�,����JK�����`&3����!h/� ��<ڙ�6,��}��\�oӈ�y�-��;�F�X�y���L����=��.p�5���?���z�C�����O�d^$�qBӀy������sMH��3ڄy�@SG0|��!v�%��D�Y)�h�W�[�����[ꗉ��3�)Ge�#y�Xrnm�do+2;,�DȈl�WD�0�v�˵����C�6��j��0�L}�Qhҧ����d\#J,F��`ٽ�5&�Np�g��,�x>�i�
��+y�3-�8��ҹ�$�[���ô7\{��S4I�D��G��}u��	7e�ZCÓ������f30�]�γ�J8��a�=��J���_�p��gW��lbJ�}�wΈ� ��l ��"w��"���iA�8�g��wF켋�Y�ǝ�,�\v�͙�e ��?��-���^�a���v:|c�]Q4�6%�[*�<Z�B��
�׺��RE4���d(��BY��C9k�f���;*a�5��}3H�t����u�an�Y��5��^(ڲ8���=]�a�D\�I��1�t$���a��w.�kc��r�o�}�	�ðЊ��g"�*�j6�{%k�����^L�F"�z��x� ��wq��D'��M��,8�IW��w���W'�fb߈_�D
8lEO������f �s��25(U�̈́}8�8��U�v"�;/}��������7WLqo��x���B���Aŏd��Rp(��U��1��/q=r��kfF�>����<�bB��d�.���rv��`�^�Z�I�XA@��z�t��-�׮
�����bZ	�'��r���i �aT3��Z��Pnbt��,��S�*逷�06d��T��А 
�ԩ�?B
#	=��Y�A�Ź��Z����ꪮ����� V�
���� ���y'�W�V�n�>LN6��s
��MǮe���a���~`���M,w.�Q�$��L(1OD?�����E�<#�*}�B�fw%y�V�a_ck
����=K��J&L�3��AA�;���b�W�A�-j��&��n�x�L7�(<οQ'3�t����;���������.�{,[�T��	�o�9���� ���ӂ?�k*�
��$Q2�5��1,�w�k��fbAA _��o��r����Jcu�̗��0s.e�������.yR]05Y�~Ӡl;9(*q�YR�xF�ݲoyPQ1�]�4�V�A��>�ز�:ٮ������R�ZE�8�C�(�g@%\֨jzB�7u��p����:�������t���1o��S�|W'���{ʪ��@K�/�P���"6��\�����g<�}>ApW2�^]q�A<�O�Sd���^�R1B���-[�/�Rh��n-���F�|��⩽� 1�%u-˻,K���ìt)��|	O��^�t�;`e�_�\����yc���I��<)��˄��9٤�a��~irh���|&����1*qEWo{����s|���cM�U�
�"|n�7��i��fO�<7�K)��_O=�U�W�cc��Rc�H��|p!˨P��KD���8��_�t�_�+S�tcbљ#sP��7�O� ��:�x^��s��i��G�è��~��
��$˰��<.rW�V��Fa*�|S#@��֙j��4N�cG�x�,�_/f9s��H��������ܱ���RL�e�ĝ4kF���d��.�hUu ��ه����M�@Q2;�M�a��v��{�ԟ0�m!-�U����y�Xw����j�2/ �����o���y~��@==�9�I��q L�d9�����E��!�����п��y.>FB0M�giN�.p��hn����=6*|Ncd[ʁ���6ua�o��/3�'JVWe8�����#t�x�����+9+�|�a*y�ĄB�����IY|[ه �U=zh/�gZ��vda�]Z<<���rN4^�,�D4R4��!ecC�	��.WS�80�P�I
��.��#ٔ0~f� :��mQ8�S�D��d4x3��s}���[.klEhw�d�y�t�O�����	q �m&��^.0�����ϗ�<�&�v�b����vE�)�v��{V�J�ֱXO���f}����ޱ��S���ۧ񜶈(\D,'��=�l�3PR�xB��H�_��U��?��ϔ�>&+�p�3<����=L��:��w\(�t��:/���򄓯�Y������z�+j��+���J���!����Y|�a�-��,��u0p�y|,�&�G��8�kD� �Wn=M6_p*2U`U�ľ���OBMvG���C098�vz�v�I��!�p���Gff���~/=5u��i�p��[�~��$������Pu,�D�],/5�}L�zǋ���;�G�J��3'��ۿQEl3�Z&Fue��#�P-��i�l�X��D�����~u�}�8���X;uo�3�y��kǧ�q�x-4jG~O�����X&� ۟�������zں�`!d]�i�+h'��q�|���fe���eЉ�ke��x�Ո����t���s���ɷ�!��ѤyH��g���~���-� D=��Bڒ5.^#Ϛ�ɦ���4R'ŴP������{9�Fh[D��K��(Q�B��X��]��z� #X�妐�OL�H1]_���u��"���4y��G tC�m#��������i�~ɞ�X�A!�ˇCD���ZO�q�w��Ff���5�{�d�Y`{���Y��g����g��� �wދ"g�[cP\j�-�ok��j nr�B�Ӹ`��$��� %1O��証7+5/l�C8P�x���h��|��R[B!������P
�G�baU(�nQ�;G�:Nq�n
��7u�dG^�刓��o}l�t@W����A���[*�V	� �C��To�ӆ�{gE�iO`C\����.4k��ƚG�����e����	�CBL�9��V���$�" !�ml�����įY]_�K�M�@K$��G��L��Q""��UL�0��ʀ]<'�pі|
���� 
�ć��:l%-w�D!���,h�Z�`BX�$���f!���r.����%}�`/��`�:!g��5� ބ���3qtP��W9Ia�~�|g0�-� ��m�H?~V�����=\+S_EF���� A}��8̡�߆���o�\
Õ��o����E�.�A=�׸c��?b�Ǌ��@�x	F�З�������Xa$T�L`E�H@+�o����'0��C\��"�[�Ѐ3���*{��i�����,r��о�2|b��qNp����`�7��	jTl�z0[�:�iT���P�a��7uK9��h �����i�/C��
Ǒ��̋KJ��UbgT�'+��+@4�7�pȕ��b�?5g�d�vSa���Kcv���W�"�15K��G0r�AY��7��p7���0��v+��$fq�V�l��wt3��0
�,�Nތν?�#���*oĦ
��hEz�B�ZP>�x݉������+;��VZ�/��R��h��3:� e��!C|��3���{� 3���~����wAW�>����}�8W��U��X`��%�l�����t@O���ƶ�|�\�[+G	�	�P6�^�r$�|d��^���{jDPS81�B�dgJ�A�DlmR��.ԣ���72�{S��F���j��ooE���߮_�p��@wi9�Kjb�����$�c>���L�Ʈ�����i�8c��P�Dk�Վ�����:�+�I��xy�$J�
9��������V#V�"J񋏕�DYityz�?{���8�3Vs���`�8v#r�%x<��\���p#\s���@n0O�&�3T���R�o,�NCN�l��(�G�ñ��/F�E1�e�ð/�^�F��e�þ�8�m�X��x_�T՚�	0��\�W��펾콻�\'�2���_U�&4�R��Nx	WR�*�c��C<���������p�W�B��Ow�fI�L�F�#�l�눘��@Q'A#i����2���T�Lcm8y�z;Yw\T�K�������n},�t�B^a���J���7�X�j�(��8�˙�Ǿ�pW	E}R8�f.��#!���<�s+E{����#�UU��|���	�'��`�t�n��p]p����k�b&�~{к��073�<�M��nӘ@R�������/F�Wg��0��{�_�������ځ��gIAꤛkz��	J_�09�Z$�2�5d}�ZQ����J(��UE��qKEI�L?!8�H�z\br��2�����;.j�b>M�n!�{���i��x���k�z4򔩶�p@3���
�YZ��g����_����%�}�B�?��M����[`�٦��8��]���:�0��a3��OϿ`[��axw ��_G�z;7'*}Y^��)Fce23.���.��W�L����z�Bs�����f䄞Q��
I3��H�E+c1@�� WL_��V����]~	'9�~���|H�Y3լu�yR�P�bTs�����R�f�}��{���7������j����	g�ϷF��w�	O���]�g������R����Ss��L����1P=⽽D�D!�z;Q���d>�g���&����?�42-iQ e<L&!Y�6p����!N��
aXz3%NFPJ}L�(�|mtm�`8�K�1,�8� �zg�H�]��O�E@��X� �U���T��5����Ȩ��ń7$}g���ܟ�a/x�∨sYT�ks��2`�?v����/���S>֮nޣga(#�m��������Ӛ`��-Ǩ��0���<�����h�$w��gJ�ũ�ҷİ~vӷy4�v.)��V:��TR�Io]n�B�~���×��n �g�`h7�~cd���ϪS�&:�敉Z�L�g	��j�3��`E�-L�m&�Z�%3�>e���f��ED|pq�i~��PL�o>r�1�8�ԭ|h 6`��Re�n��!��9��f-wS^�+��g��<�i��<;[���?���X5�>����ꃁVek��S^u鐁~�����Ȩ�T��C��Ȝ��k�Mr<;u�D��v4�:I|�6?V1T��2U�Z(�dzx��\!�w�+	��Q'Z��e�=�	�^��|t�<���~�[�$�|s[6)%�K�i��{�_z�x0�|�v�aI��>�7���-eՊY(n�N�Q6�.M�H3��1)㪆U��W���X����֫Ï֠��f��m�@6K��_��	v��B�l�>�wM)'�S#��iT�	֮�����nH@u�G�>KIB��_L�k�ȝ��O�V؋�?#���t�
��?��U�]�3ri}��$������4�3�:�b2�o
��<��s%ZS��\YW�DlD��U9i�OYS�g�-��L{#O(q��3��h�y���G�~�tBR�0]�1}4Fc�5bXm����%0|�k��7:��Ƨl�F�M�����p���Y�.��Xo���^�\��ut^G���vٕ�ݮne���;�Vc��p�!�eԀ2}���IS�6�����WrО�0�H�5|z����.q���Z�����L)8���i+����/��㎾���H#�nh�qX�R�+aa"v��.��>\W�"��?� �>a��Ü!&/Yu��>Ȅמ���
H��hR���i�
(�V��钺?�d�~�e~6IVߤ%�rψr]����o���)9�V��A�ѯ�8���}j�K� �Ԛ����V���#�Ȏ���@�h���-=hK:�y-A΢=�,#��;%|�N�ۂ�F�8j^�У3�_Hu��l�����M���źI�C��[+�v���:�x�X�
���������u�H��W'2���j-���s�vRc��X�׀,����O�Ն�]2��6jUj���]Ľ����9���i7�E�OH{p�Sʱ�K�رS������i� "��̵EGd.,W�h�XNlAf���Ɉ��iv�2���N[��|L����0�B��=���_�{49O�ߝ9��
wX���݀�8秙�[��6!p>�`o"���:w�|!�K�PR(��j}["������Oxp�,�8�Ɍ��*�f���	-%բ��۬�"��>��ӼM[B�\�`��*��g̉�
�z��ş��}��8AN����*lZ|��f�>��++�Z싯t1�h5�~�-��4ۻ/]?ah�/8�����@�q;�����/+�rD3 AB_��ڳQ��P� �F�O���Pu'Y���y�嵪s�=���GؿG7҈�`)�VQ� �V���(:[/ܹTx�L�T�a�d~�(_"��w�s�՘��(7�������@+�`�@�9�F|oڕ5G����mJv��n�؍l��P��y��J��R���O�l����࿒�RY��$�V�j��I�C2��_�S�U[�������uo���^�����:l�����)I�k?�f�-JkC9]'Qs���[X�LU�#�bc�}}��{9
�M�I�yN+���� ى��J?<=|א+�y�Ǘ��!%�TL��F]�a%h�>�f+���m�r��{�d��t�D�����?cQ���{���v�^��;*��z�p��x�H�SL�n��J1L�6�����>�x&��nG�b������>�V,���{�O;�Zq��R��ڿ5�/��$��}���?�J�/�ц�T�WIy�0cМw��j�̜��_���T���>��C0���E $B��`gI����h-Ֆ&�]D�X��]��}��D��>хDkye7*J�׊�O��;��w#F�L�?vo�P-@*+�˽,!�E?���m��s���)ӓ�.+�%��P<��;/��J�z�V?��8v�4��a��rd�~ E�@�B�G餗�F4_%�Ժ�*%�O�x;�W(�_e�Q��
��iW��I%rG�n���J�x�K�Ӡ.>b��~�ub�҅p��:\PB �T�C�&�p�y�HQ�{�������Nh�pnx�i�AD���,kD�m�w'��"�J:������Qj�j����W
��,��8�y<ց���H�fSF�$�{X�Տ�J�k��	~���l4�jK�����q ��5�<��,�+<��=`�-ߧ�Lgú����/��WOh'#�*L���9��n�t�L�`P&Z�Ȣ�1���.�qE�܃=;X� O(�CW��-��Cľ�\��[E����r�m��Z�KD�Q&*�� ��.£�qC�k*N �t|w��g��Wxʅ���?�E���b�g �<2w4ҶB�6!�d:�GѰR �����։��>=ƼD�P~[�٣�s��7����5�ל��+�b <y�YdS��MmO���.��t�E���߹�6�1������q�l�_��~R��>A@[	�tv+*b�EU)Զ��M`\��f�N�G��a��V0��.٭��e5۾��Q����Ӗ�=�.�@�����D���y+g�jט����Z�zX)�w��S`�ejT]^@P�uLm��KIZ
}�Z���@T���D8�:u��𑥝�f��8Ϥ������t��6�kt�3(qߛhpN��}i0��4.a�m�c%�6��f��^{��p����͚��/Ga&���3�D��J���qm��cbС�Q�I�)�z�����lZ�9����Wj��sW�s��;�auX"=^�m_) �j��V6G��`���R�#�~�{�с"�dQ~V�0q
��r��.�S�Zdt&��d	�T��ֆ�8�p��b9a#
�&kYx7�n&�1�&��_��D�,�a.�|��۱&/�����e�� =�4)���?!:�뿵�Xp݁y�o�ꖝ5����U���(�-��i�_"��>u�@
���_�r�܍�bg��]���LC��C*vA��нT".oxa4
[�xݓ����3��;N�ڲv�e�+ա�|���k{Կ�3�^U֛~	G!E�����F�9s��ZJ�|�Y�5�ߤ��t�}���A��W�gR ����e�Շ���q��=���h��?��v{�,���8�T�#�J-����jq�<Tcd\��9��r�4Q�(17�տ6:Z�o�6]̏�z���Yf�"~}�[ |(��1�$�p~�n�;�G~���m������Tq��&�=IN����(����?�(��i�'uU���9���ϑ��}zع���Zy��Z��P�ug,N�1���!�{~x�6Ug���O�?�W!v��9��k�=Ya/<�A*@�x����w�|Peav�Í$`e#��#'�ϥ��L��e�"����
��q�V�%Oŉ��do�z�jeڧ!�d��.��ɏh��C��k��;"0�&5zq�φ�pSlp�����q����F�U�a/�H� ��M�^����b�T_<z��-��/�V���J:�$A�a(:#��/<k�$���R�[��Ʈ��sg��Nld|VT����t1�+�qQ(h��<�HN��[F}º�le�9�l�ʜ���920m�!�o����eA��X�'��
�����g��ΰ��O8��ӞZ�1gp�P]7���®���`?ZV���4��"뻏0ŠG�;�Q#�!�~#9n�Jm�?�X�G�i��̳IR���R�1T�A�yf�8T�o�n~~ބ��X�^�%5Z̮-���gf��uͥ�)�x��@����5��f�3�D��]���ت�l�0������4����5N��]k`��-8VGc�IL輍j��Ũ˾����u�����l���0��C}C���᧺�� P�ѰA�8�TY2��>a6��p@Č=��%��v�S��/
�'�S�{Ѓ��J�ؿ������, ��m_�&U3}���4�5�M�ְp�K+�S�r�C�v���b�@Y
��ǋ�!�9U	�Pv�D��$p�G~������ǉ.�_�f�#��D���Q،s\��@cs�岫/�?$4��O�C�Ѽ�dKW#��w�xD׫�Ձܞ��V>�i�;V�+��ǣ~h�/���Ĩ���Ǖ���F�̳h��A�����@C���T��/VNc��/3{����]�H�~[g��D���X�"x��+�)�*�ש��d��-#aˠ~�*p=R[�ԥ,����2��sG�Q�4�*Yy�=�R��Q?6�@;�4-��g�s�5��H6{�
ov�5�1�M�\^��*1T���!
w��?_XD��E�l�9�o���Gng�Cq[�%(f @]�VcQ�EMvՊ�z�щH�)W�#�L=�D�t�_�_���v2�bM\�O�D����DL�~_���m�P��4��ex�Zv/�`e�~�"|:��	.�lG��0�'hp��zC��0�����4�`���>��rй�p�CoS�}Zn1f-� ��3��9ү��2���t�4wx��������-h>����"�!4����ݷ�y̪�����j�,�>�6����M�2!H7�W�z+��WՂ����M;B�<�P��G�$�nt^M��f�G�H ��')}�?Έ��FAt�{�Q��vO�Yn4ԍ
��_n53�*Ǟ�x!�1�>d�$��ᐓ �-FA�ePOu�:�Y�{+��/���:Y�:<��/�ސ�h�����a�2���?�3-�\�N[JC��:c��[���,��L&3�.
f'2lӲh��jlU+jsd�r�8YQ��s���!,�D&^)�4PY6+j�X.xɛ�{a6^_���t����~gz`+��V��a�`���A]�B�.�q�|����� gr�Y�K~U,n(�[�Z�� ���]�[`Ikj�s$��C+����37���uɀ�ԃ�{�w��S�ǅ��hW����Y	H���إfn	~����荊oEq���p,��ia�7(RP��/�҄=~�	����~��VN�Y|�^EK���e�vn�8�e��F'���Bx�r7O���8�cD
$_ ����N��㚠7���@�g{�j_�t��R��D �0)���ߘ+ϥw��΁8��7׵�8����6E�q���T#=q�%�ϑd�!��z���of����'�3��J!��=
G�[n�b�ṭ��y��\qn���i��1H	���x��� �,�Q[� g�5�M��fP��n�)��dB2�%�>CM���Q�Lrl��AJ�z����1J�m�IsN�g����W`�h�mo���=�8)2N3��Ӫ6�w��ǫ�K���M�uFp��"�^�ŲQU��#�s���+TM;���#��t�nx���&/2|��=D#��KH��ņ�/H_������ǥ�8)�7���RU�l�:���?����D�3(7�h�
�q��ӎ�_(�\R1P^d�o�A�|��M�N���U欉ڈQ��U�Z��kL�0�v�ּ�� ��F9�[��>�
�4���5�D���xgsPrD��y�� ̬c[{ڸ�qe>+�����e/��&x�+	��Q»�v�[x!b�����"�`�*^� %�j{%�[ȟ��w�-I���}��C}�Ҽ������<k�W t�$r�nK�`�?��@��ʻ`��u�tLM����j��ü@W4)�E6�	�qb�+��7s�}���ʱ.6$�y8Y[��|$����`� ;e�Ə���He�#����5Z3Pɺ븻d��\���~�'Tyd��H�"�^�L/����l�且L#P����h8
��������ߍm���&"o� p3���u��`����.q2(�f_9�o�ͪ�Y��W�� ��]�����L=
Ki�0	�Y�����n!w�Bz�R�B'	S��TD�$������Y����wg'���bki��¨D�ˎ���䣶�ю$]���wDzt��-C��t�C�n5��w�����9��m$g� ����悃�1�vJ�]�`0p��Z�`�TR}�'~H�&�q����9eg.�j�2�=|vYEz�n,;l_�kq���&f}�I\�X*��T�'m=�S���#l���^H�?H}�+�YZ�\϶��<r*�&D���ft�	 �|*�݇,9#�Hz���lCz�L�0�����^�fq���ݝ�1���8�_p۾�,2A�Z(���0 V�F
f��[Ά]☽���E�e�dʕ���$/����60�%Ō�[؅�ˆ����`Ѓ*��%Z�V�H�'Cٹf�ŗQk��-{��m'K���<���=���іҩ��{6���B���T�͌m�w C7��@q�V}��j��"Q��:X*$@�`�]a
s�ԟ�eg�#r΢����.:�n#,{��nV�<�1�-+[*��|Ӏ���AI����[�_���@~D�4
G�4����4ޏQK@���E�.��m*�� �eo"������_%�[%f\��Ā�q:��1�-������kZ��<'Alۼ��o�A���熱/�!��aJ�K��<����?�y���LB��=�z���*]]<�6�|AH9���=�5s�B9�%Uqw�{<�<�댜U�\��#4&<3��^�B��� �έΤ6f�ƨ=��1��QjS��o��-y<��&6^��᜽9a�T���:�j��G:ʸ;Mo���߈�-Z����z�%�m�+�/R�/!،�Fr����7v��uY�N��n�H8NQ9�����w�czWt�G'��{����^��ó�'Ofd���N]�ȵ��xw�w���r���`v�ꆹ�'�u��6<�Z��ޅ�gڡ��4p��	�Ghbg'�Z���ـB���c�g�J�97G������bc�nӰZ��L��_)���(� ��l�0�Z��a����G��Ϻ�˯�$�/����#�ս�^�Y��70�����re*��N���)T���*N�|MZ�yd����/�'��;�����#�3݆Ƌ�`w��y:H9���8>�F�G�"Ŵ�o& V�Tv#f��5����)4Z-�ѥ1��m]>S`|0�6�����jܓw����P�^�h��N�XХ�|��%O�cW�����'_��V1zGeM�R�N�KH��R؅(����Q��lQ�>iO@��(Wc>����O0� �G#ĳ�Z$o�3�������������� ���]� "���52��pƗ�l(豗j��D�D��0��֏�s�f�:�,5I�>��q��Q��3����&�ps4��~f�T�,<ɉ8F{s�M]����#�~�����rGN�gL�3�n�)L������4f�ye'�Y����6j��9�<��3�p�b��6+!U�	�_�9-��ш6Wɖ�t��	�:���k#�S��jk��CPk;i�G�!Q<�S_�	�������˓��hB��lY?uNT<�������_~���@�,I���F�m�!%�w�#�r�7|!��@xW��~rI����+"sg��c׾�:g�Q�G��a���>A����qw����[8�� ��v�}Ba?�J�s\���@�|�n�JlV��= �s1�+ g����:QK�0��s�jSz�I�)4�����`�(!������C�3Zh��a�5��Qu_�W�k���d�����YvnuI|ɀ`��3��`2�)�/�6�|��0v�
o&]{:�m �=��&�ҚU��J�"��	���)bf@��X��Y�O}z$[�ճ�}~���)c����u������p:D�� �4a2�_	�Ɇ��f��>��.R4�<H��goq�Dg��Ǜ����s�%Y�.�R�:l+�<0�-`E{��k(#A��i��1?G�r}���e\;"���Ȍ�V^�ݜ$��#�(�e�I��%{LP���7~�|�����j�0�8�=rF২���k�l�-�К���y�f��)4�X�4m[0?l(N����rn(y�������n�j`��z� 0\���lJgO����Ȉ	�ū��^߈�4U�w�	�gJV�6�pNs2L)��bZ�����'"QZuIx��l���z�,�ےL��@�nJ�T����`f״0����g��y����Q�ן,2Ow(L"N ���MO���ZllJU�jEC���1�+t���O��'��W�6���.�L��2[��S��c���h�]�+M�n�����N\%'�/�����=�&�(�V��l��f]{�=^1���j�h�-�`<ӱ��.�����r*�k�d�e���η�=wa�~������8���q��]�Y~� T��z|��1�#��-�	��#�P�u��ׂe���]O"F�Z����q;]����F�R[]g���^�ۻ��؍#�@�1*�>H>b�H`>?��
!(�АOff�h��:�ͳu��w"�̽�}"�y��,0NC`sG��p�����l�vƞ�
�ˮk�s
�X��f�p�W�����	0��Ȅ�)����w��N�/P������Ǧy��O@h�r@��?��ן{eި���)���/*	�j��]��Ͷ�y�5�K�z>?c�Ƃ9��U�]��A�=+7皮�RT��'��s��i�yj�����3�1�(���cׁi��{χ����3�^�RG��%W���o�g@1��X�:����J+B����t�|2I�����X�*�䥦О)��%�������:�\?���q�$=��������~.��E>�o%�hM}���`�@�M"�`xbE�}�D�H��F�T<uy?��1��l�5��q�Z�K1O=��G�dۢ�v<�Λg�A��Q$�_����Xm���򈣆�x�*�&}�����
X_t���)�9(Og������R�_U(x��ak�|����[
*���2֩͡������4��P
�%�����ȏou�e��a7>�>J�|��xB��0�@��e�hY(���l[�ʁvڲ����\ǢWoqb��lJ�˽�Y]\X�R�3{x�c��pZ������[g��V�w[o�̟��Kj�M^X���z����y�}v���^�L�������ƑD�G傶D�i��5�@(M�&����̨]��`����W�Sɀ�Za0�i��.��3f��^I8 ���j�r/m���l�=o6�1p���3h~�^����N@$��� b�%g���T��H��1�g�=gG>+�>sz�IRH9/?�1�dM:�A+,KJ��oe�-I+W_��3��4�u�M�� �y��#K�lQ2r�7p2�21py,V�Z^�bzt�����ʓZ�f��n��,�ފ��W ���j��[׉��G�
oG��;��u�z)������Р��Z�	6�m��MÄX�VK�z��|��ݝ?�PbQ���6�v\vk�dH+x�9��z��n$����&��*'Yi����"6�y�w|^P���b&sL��r��́�4�T�s/�Y7UIǴ�!��?�i��a��r�_6��cd'wW(���ňOO����#Za�3���E��V��iR~��~a���o��{|��UVW�ij��,��3ύ���M�ߙ�L~�z�糳�qliA�@z�w����Z��Q�������?��g�b8��oTiH�nt�/,6�3\A��R���2:�$��(dW���	�"��fE<HI��'���z��ucw��N����e<�h����%Ő)|��⨆h��uys�:��gĸ��gT�N�Or�p9��G�m��Ҩ��H`vls����φ�(X��nܴ�F��p��8�J�'Qo7�����\T�])���4���Ą�w!�W"�:ly�M�I�����A��zs���ec�,��u�j�?�֡X i��#�s��H7٨����M�e`,Vrq�d��vQ�`^�~��o�5���f)�D�����m3�Y�˲&��8�x_�t�.���[�7M� -�>����z�j-a\EM����D��L@�b�����,�*ܶ+����	��I/��2|z��ш���%�ՎBH�sA�5�%w9�C�s���<>��1Y^|��B"0>��D!Fk!��ABF�/��ϋ�6!Ӥ�����K\~A��E��)�z��8�ĵ*�����w�_�ɇ��ʺ�å|���i�?"hN��Jܰ��ܰR�Z	6���Ʀ�բރ�?��uu'(l'4��]>&�]\x���_�h���׮�Z��T6�a\��X*��UƑ?'7aZ2��� ���iW#�t�mN�u�$���g��hsN��$6���8O�E�4�I���R$��Pc�&ͯIy2G:�N)��$vE��������S� �D�D��^�x�]Z.��,^��j��9�\y[�/>Vr(2� �A�����'�Pµ�c �MT��hA�,%��-����Vlj9Z�Ȋ�sFo�_5J��m���B!���L���z�����$�Pb�����+8�����,"������v�n�ItkI��4G���� ճQ4U)6��.�Fmؓ�x���?)m�+��AH8%W�d�>�	(�4�S�97��;ǻ�r��j�Ruof� �7+��C�L�'�m�~�Þx(�|[�i�	�ULB֎7�n���g}8�F��i�g+|������q'g���a}������ɻ�Q�^��s� �[D�B70J��@��l�	��e�P�/G�S�����A�rm���"��grI9m7������b�e���7:{%�Ăd=���:3���h��OD]R����
�|��>uɐ�Wd�ٯ��x5��9���q��wD�*�Xj&�iBI�g4�� ��3Qg�0.���]�� ���]��v��O�)�.k��^v�!�<#9����r͡�f�����n��J[UC�<�W�G�{�x3p[E�D�?�L�3㾽��!?/���ϭh��Ωq:6o�:l(>�=y��0Q���Y]����>���h���`�IS�|�&Mj`Q�Z<MI�u�kL"�'�޹t�uC�А½	��N�$�i��M�װ�"�Y�ʓ �%�k(��f����'��"U$.W�|�Z?�qV+HP���E���R�2����.�����KG=8,ֆ�P��U(ˀ��u��[9�kzy�Zs80��ꍱQ�OTa�q��ҝX���Ύ�P�~����ca��p�`��W�D�\�`g�:kmDZIY����d�k�td'*������<�?{΋�D�V1.�	�[>�}�Kre��/`��Q-DiB��e��E���^�lyaa�%���H��ÄC��5�P&L�I��w.��H�m��y%s���`4��q�G+���Q=h�g?1��d������-�rM��}��a�Hَl��#��6�	��
��#��3u�ٷ~�/�	Z��./?��Q�W&��LN�s�[b�����;��6s��]�&1#�6��F����|P��$6ْ ƚ��XF��{��g��
����?Vz�8���n�Sa���!��׼�w��|0MW}
�LN0Y;W�9����ö���z�u�E݁K���1����a2i��Pd�@Q�����݆����&�5c�S��j�?aÏ���)�N����wD�2L����Z��a
M�sl@Ͻx���Z���q�f2��#�ݷ�D!A"�ui��|ct��^�Ɨ"�p�
\jcna�n��� ؼ7��#���{�s��H�۸ $��<��)�O���P���3���RJC&)p�����-�_}����s�nc��C5_�.��"�m�=�*�Rta�Zh�`�Y�[Xy �����ve�Q~�M��Dg��p���Ǐ���/�S��Ni�~�+�=Ĩ�� ��6d��7{}ĉ�(v��\�U:��U�$/cn%~�����ĝA�C�#�2`����s����(�����:����S/�z���j�&����g�Y�����6���&�2'�*���)�0�㸸5���@�x�+F�OB���zK�Κ �p*5����De9.Z�^(,���ϱB�^c�m3Ԝ�Q�9�`��.�mJ��r��_.���GŒ^�mh��]��� n��X���}�1񅑁`��|��w0�*^�kV	ԁN#���!65��d�[tM<�%d�C���O���@�#��Y
3ߨԟ����}n����D[�����߭���\�������րb��Y��=��׾���
R|_�ȖuY!#l�aͱ���ͥ�l8���jŹ�E�à��C�0�Կ-�/��#U���%�؞k��݀����;�(��9��p���0��h��g�O�m��5�g���L�����
��
��T.s`��a�:m�3��c�����;���C�-��x��U(I�b*�Q���dg����=�B�8- A�4WgT�-��U�"����� 3D�ș�1�]�O�a��x�r[���d�B��w�x��!ߖ��(�;bv�P�8YF�Y6���G����d$�+ƣ-���v��+ʑr��,�dUy���m4�9q�T�	�7B��QOď]+�D�H2;���ڠ�)�{�\F�c٨�ŴūTЯ��kG���Y��j)m�$&`����\j��K�6�	�@�o�8�� �Nn�^��L�刱��b�d�^]VX,F,�@�,z��E�O�ۨ�E6,����$��S�C�O��W�]�b��7��X�v�Z���G�}����?`-hƂ�м����s���}ًځHhھ��l�
2��!�JR=�_����f|=�0vxǉ�b���S��'�+믇�l��ܻf���H�m���v�t�ʕU�v#��n��]N1$���7g��� �;��	�� V�Yő��>d>��F�;���1Hg�R����|A�E�-��KȻ͍:���4x��	U�2�8k���xjW&�A�h�!B��J@-L��5:O#f�X:����`�����*����M�b��Bv�]sFզ�R;�W�,�� �j�>�����*�@<�sط���m��Hb�\5�:�ڂ{A,��DU0�g�Pw����~��>���iV�w�_�)<J�B�:]�g��z��}l�����;FF3\��O]!�g��X�K��+����Ʃ�^s܃;�0s2��\�	��U�w!�RE+��U3آ3y�ɇE�
�j� +�5�������VZ���>3��B�u�kBw�=ǆB|J�n>v����n�~�%�����^�F4���x'V�$��y���3�O�_p�@��,�뎜N�6�^.ui���E�9�Y?�!}a��d:T�fl�,0!=yu��L>Bo�#��Ǡ�C�=hM�a�A�Qz�����u:� xΞ]��hh����0o�����f����d3���F���^���6NAҵ,��wo�p"�w���S!;�����e�i�}%K�,��9iH9�z�$CE�@U�c7ܚ��ˠ�f�������S��O�b���kFSZ�qO�Y��|`�������K�3P�a���GE��Iה����{ s�5��ia�]89
M�h�E��i���j���w��"����k� �w�GJ�]:�}S2��i9����#(�mS؁���s��|�	OR�"����(�CF������Qo�]S��-��tk��v׃�Ĩ���6��+Ou�Bb��Yb
�?jf�.S=����Z������Φ�����"�Gu ��4�-G	i
�4�^J�~�+-)SE@�A�T��.2�e��
47Y�F{9G"��߲���?[q����EvV1��k��^Qu�)��2�v�%BP�������M�}�b�R�ю0b[���lm�Cd�~�7I.;B;��Pw�
��ɪ���#�Id�j�]�?���,�p�L��a��
H��!>����y��#�C)8��߲���9}HF�r��}ˏ �eQ�u�^�m�/ĵ�z�,��|�ʂȭ}'���RH��u�5�@�����D�
�A��������0U��VfD��$��LK��W��z�����9��c�dd��Cl0�F�:�N�4g�k�d��_�}Q�fO ����$�W���xV�.]7c��&lL��}�d������� �R���#�eo��qO�h�G�z�>�X@���^��߅�H˗�}�:a%�o� ��F#�C�K��=���e*�e��q�z�1�� ���x.���ubjm#�����֙����b�,�CF]�������l�r��Z�0]��|��,@�='B`��
�����g�þ��ë�LVf�C����<�9�^o��M�-�Qcג�S�sxչ�H_����[�<��w)o-b����N
�X�N��T~Fn"cM)�s׍"~���;寛�-�2��)Rv��D�>-��%�ѻ�oP��T��A���KXB���I��0ݵ�0c�:(^b�kӻ^��Ů���,�}�2���E +p�𹩠I�!�4���a���,.�M������;�b�RAvҊ��'�G�����փT̾��o	�IDE����z8&���?��w��`��(��U���cf6P���<j��/��UF�ʀk�Xx�� �<�����+@��7�1 l��,Q�!c��H��=�w;�Jw~��r�B�����x���"ȗr�����nH��##�W
0�h�
�h����ɡ�*����>P�>\����𿔥S8)����$`��R
٫�&��<�F��~��ɈʐV4Ѧ�p6�g��i]�$�i3�w�b[_�ӡ��<�������̓"Y�e;�������.l�.��~���*��?�?2��-M�Z˫���A���Q͑dB�
^lTxv1h��z�=1���Ε���#6��UYQ7ǧu�����R��9�ڏ�:�l��ܜ��6jS٨]j{��E����|�x2&��?U�k�	���a�4�������g��}c�=VAo�� #�%�swl�x�}+".S%�OK�
Mf��ߜ�QR�F#X����f���SX���z�F"~�r�5�3�|�;1M1�/e7����T�=)��M�\����\��|�l�[A�	�;�}��s *��ql��x���/1�䔢qNO�N���)\��9�}9OĞ%�{���DI(�]�u+�� ��4���:M�G��؎DS?z�R�Z��?8���|�rJ���0�-�G�?JT���Sqhw�du�9w�&k�R��xU�Q�6O��dl��qt���' ���;j�!�p����,�{�	�/�?��[@��]�j�s�v"�����Ԭ���>`���v��N(�@��7�6��Q�)�ApՒ6��qm[�ɰ��>u#�HV�Қ���	��e|�o �?�Otmddj��(AN-���E��o�bCj <,8�C�q
>Ta����[O
�����N����t�붼�T;��0٢���FKS0e���r�e1�c�m��r>R]����9�?qs�T��N�S/��.�^|����i�a����^2.�>ţ��.HAo���g-�A����0��Ti�1��6\ʦ���;U��1�6o1U54~�Q�iq��߆s!��`{��]�bqC����<N�Sm�(}j6H� qts����]w�,Δ����)�/ȳo�oQ��w��N�i��S��������'�8��m���/}�L`�ˢ\mYhǚ{2��w��ͻc`��n�.Ø�n��_�ε�<s���NN�2e�͍���	�5���Q[`{���!�,�����	��?��u��9n�g�G�k
v�=s�3U���j��d���/'�r�? ��i*�_�swر�H�d�cr��Ȯ����f_�@i�V��9�I�Zăl��������Ќ3 tŮ�~ճPX��Rݤ.��X���4�����#�s�\)�E.�0����o�O��,|
��Ԙx���1
*u<�ƦE�t����$f�3?M�'��\��7׹���T�
�70t_���O�rY��R`K�.�M9�s��!L/��ɫ:i�0�=#\�o�W�����@D�R��5h,�3����^Nt�I�ܾ��ݮw&�0q�.�����	��E`�v������.���&�x=�~�:�D�o�P�H?i��ߞ����f�Y�3����?9�E�ӧQ_�P�*��m��X��E��������b�N�28~Q;}D����B㐃���6��ܩ�T�C)u���z��	Y8<����r�T��e��K� ��
]�9��?ഺ�䰼ˬ7��B6�r���3H�-<�Y	fb�z�O�@�`����<������
KUFI|�;u��M�}�ޅM�fQ��B�}�s�kΟ`�������8�A����ְ�u`�8�q��`��g�	QZ��4l�N�����5�*�����(�B�9孳�����D�əH��ɃJE��d[��{;n#&�B�((����>�$  3�{����%%ɿ��e�.�R���O?���o��qܽ;n��p�E���3L��#�S�Ly�d]�f�T&�-p������<���L`v��cЍ�S�L��vr�3�%�}��h��Ɏ K[��Z���"*s��gc?�+�$��&�,�	&������m�@��6r�z��X���ؠDj�9�G�T0r�<1 ���K##iM�͸%i�M����t���f#�0�I���S�[�T-�.(h|��0t���-B�B2!�&6㱼��W��������)h���lĵn�mb�a3f�'@�a��>�G�Z#��|�z4m�V;M���_B`�a��: �U�ftw8*a���S�gu$Ň���$n��|S�Όa�L(9G9��0j��U]�"�m����X�M7�|��ޜ�����5�;ʇˍ��Oǣ��T\��@�^�g:�a*J���mW`��ϐq��ƙ�J����P�p�v>L]e5���هN"��¨1��@��'� ��e
q_Y�Zi�<3%u+Yz��SrZy#��i;���s�b�v����_�����O��7HU-�]L�z="� l�?��>�.��iڝޒ`3�*�d��~��|��1�$yf��=k�*0�WP��,����u_��?&rV`�����|f
�3�'rLݎZK��+����:l.hM|�I:6�[�#����>��χ5$��OG*�d�Ӥ�KB7޵ZR+O�r�N	T��	?�?򵐘�C$=��-�,'�����;�R�tQ��~�ڜIt�h�m��l����Êj���-�cvH�g���/6�T��e/���= ���G��$��������U���� ��3z��ޖ��T�㱀�ʂ��k�Ĵ����χ8%����5�]2�Q:��{�S�cJ]�h>Քmgx�ǳV�t�╡��6���UZS�r�ۃ�?�*��hei!�Ƌ�a�@�d�b4��J{��J����FY���+C���~-)M�|=�2z: j٨�0�N��<�`L�ݛ�f ��@�ŢE:�a���{���=;DF`k朢��y�3g�}�7����8������R{
0E-6>�z��թ�f��3�,n���Y!��C^�<����I�6�.P�m��Ά���w�9�B!�n�a
�.��9��C��Z}�u�	�,���<�-	z�7��}�t���>���I��Mgp��=�����AY��V#}{\�,gtɜ�H�
�(�]T��Xʆ���O8�D/���v�2q��=]	���š�H�e�xG�L�<�T�]���&��u+�{W:�cfP&c���ɪ$Xy�,��D@��3%�sD���#@8��	��ԓ��!�0�n���O��fEz~ξ4hL�o��3z^�&c�1�]A�����%�oj��O�}鞙f�  ��b"5xy�]��R��d��)���,����Fx3���u\&*[�+u�)���4����u�w�6;�ηs{F̡��	y�Ȃؗ����F*�F����j̮V[��S�EW�m굼�[՗�B�c?o�Sc[���|{�W���,�-��e���aL䷚�JN��Gy����V���x@���^6�P��_u���U>�Z�Ԛ2���c̒<X��d��S���ְ�b�bU.������#om��X�vڇ4�$j �~8,X>V��x�����*��4���!�N�! ֈ>�%��}�q���������sJuR��-I�SJ~�["F ��{�g�pT��}V$q��o?0��j�`'��a���p8r�/��%�!8��x8��_D{p/7ș$y���MOƱ�U����#2�2W�Z�?F���4cv`�I�
w�B8h�� �|�!��קn�t�q2�u��}34�`�/;��nx\5�kf2�b���~������l2:>��n�yLP$��o��j��#�F*�f�N���x�;
-���R��
; ��8�7�:z���,2O��Pձ��/���[��noQ1�u�7Kk1�ɘ��\@�������bH]
� ��e7�9H���yK�����>�V��j'K��n�="�U<l+&-'���î�
Z�'4�jj���PG�?�ڵ	c�p����q�.�!�cˬ G��h�j\��`ȁ�p��2��ɠ$�M6ݏ�l�����X9Y�m�q��\� �_ɚ�n&6�"Y�s�/5�	�"��<1B�Z���F�D:����a������j�i;���bI���m�eM��`�&ǃ6���;e���G��kⰥU*����]�4�I��5,1�N=\�>	�K����}�c���L�/E���Sf��A�k�_��$���i+�y����C�^%�5��D����؋EZ�ؠ~��T0�����Ҙ���AC�����PSql�A�F*��q#LiS�x@��-�" _�C/�qP�됞�R(2�+�1��R�ֹ%8��o�ZVn(�Awvֶ�T����r��
8h\��+�*� �`^>$��Dj��N;��'�(Υb��9ȅ}����@����J���BB�ث�ܿ�6:zsT���&�=�)���ˋ�9����%���_�I,�d���j�*�}�X�BHgBB�$H?H68=#�X�ҭ��+י�wZ�J�$��iެ-��x�ْl^��D����F�����h��U�1;D���l�����2/B�e�ޖL9��W��iD�ǹ)ʂ�F���=D��2�{[�͖FwO�uڎDC�� P	�{=�5ql�)���0J�����,޸� ��QI]��������o�j��"Y��K�j0��]�-�o�HGp�G�vXB�!Ŷ��&��-Z�(�f!>�B�g#Ј�{�׊��'z.���}�wL�]� ���Z�9��|M}]�����7a�Q��yO��^�Q,�Wg�+Z�F��qZ����b�<.Q���]}�����o��͎=a!�
Ԁ�5������:��sz��Ƿ�$���(��l\�Y��]Z��<�:�,�� �A����!w��NU�������~����W��vf�q�q+�(�<P`���_����mp���G�iIm:��gg�i��o�fC`O��acA�H�ۜ^M�Tr�;�Ԥ�kmE:bɝ���c�}�����:w�;9Nr�.
���'r��t����Ua�`) �)��XD���H�<��,a��׈�ލUD�'�����	����Nm�$}���+s��g��A lg�Ut�Xg��@x��L}4P���Dz~P!��H�ڛ�џ�EA����%,0�l�X������Fcһ��a����ᒖn�,פ� ��ω'��}~�4�t��㞺�6���Е��[nW�&VW?�&&XZ*�"�?�Ű�틘��<�1��H�.�G�W���$Yi�I4b�_��	��0�� j�{$6z�f�ϵ�4[��I�u`�:���(z������;(��{x�SS�U@�����Ԅ���d��tɷn�ހ�<#����7x�����#~�T�3,$^�A�+;[�o6gܝ~��teR¹Q����f�DY��k8��&��6�zW[6��	�Q�'ɔ�Pq4�V��Æ�[�a���ʢ��ր�13��jJ.�.}��Q�Ď���aE�=6H	����J@���}ݶ�P�0��m�gE�p�K���g�Q�b�&=f�qD���B����% ���f�)����Kx�����������a1
�����1���ŝi��X�9�"�LzB�I6�� �wU�0ӊ�Y����sfZ��W�/��;���i��W?r��ӟ"�1�\)J�Sq��o?}+��h���7���Cъ���N�*�c���ua��g�GSG�Gmd�;���=n���)��2(o�+?�aoe�g���[�#
k�f2� ��I'���ɔ�"�=8lq�Hb��A$mrt�l�Lp9.{!�j���,��嘊�` aR��!;d�9; ��JW� �����a�(k�½C,[��8M����I��Bυj|���"�ȿ���L�C�/᷌��
���m�Ur)l��n�PQ���T����mۙ�q�D��ű
R�~B�m����|3f�������L�\F�I��/�{��w��f.M�g�.����gEd��=?w��-\GY@��	s��rޥJ�����BG�th1m-�hZO����D��~�uY���[1~"�$��C��(s�}$�~��������J>+��@�8��.ݙ��<\J�4n`c^������5���ŀ<O���h|@s=ғ#�i=K|��8��������s3�C�χ������+�+��Z2$=��7;�g�9��w|���/#���v��{ʀ����F��ܽ�~Y���6�BdJ&j���l{��vWw���Ѿ:;|����S {�$��I�F^�~�-���
�'���t��nFɗh���o�*ZU�Li�5a�6T�u��E�8����Z!:�k|��W��}%$nY��j�`�p�/F�a4Qk8 ��p��x��r8�v���cU���rEY�)���`��%���]Х'e�;���g� ;T���u+�{�sZv���*To��
�Y�<�v0������*��mv��tżĸ��F�y����x�-Py��#L�����jE���g+����%4�qY��b�k����C �?K�&2�s5�ӛ� �m��*���Q�����yl��f�M��"�T=^?n�~M��ߒ�����#f˝`��r2{:�'cU#8	�� ̨|�ަ����)w��g�[�<Q�1��1SxnQ
�� v�z�._	�3�g�M��o���������:8@ c�nC�d+�ڲ1�b�S��Xd�*�ǝ�M�ۻ"KΨz~�G���s��͹d&�,��;B��k�>/�B}�F��UڀŁ���ZEo��e��Sƺs��u�,h�nh�'��S��Z�V�ۄ�<��Q�p�|��7ô�W}HkɝGn�y>"�^�������f�F�+�������U#[�,�h4T
�~��^}�J�*�NQ
�aǝ�a���u����}��d�!�I�ΐiD}��g|�)����B�J��^��82v`'��%��b�����@�����"��x@�U��'�|�����2�N�9��q'��'}p<���15>�s���b�A��<_Qy?�!��"�}��	�"��7���������N�:���DW����:3b����l�Mb�7'5fIt���É��?�ѳ��{���n�ýk�U&�h�cV;O�(�M������ꟾ5��CҢ�>GG�'�Ny^/3��
�q!�;��{���Y&��b"�C=n)���3l�Q��T���/����]O� �j p��>��h(�,��M_��?~�ټ04A����{��55���;J��%y�f�����ʑ!�.+��b(��j!L�}�@���0���k��(rPΝa�����v}�s��6di��U2&�\�/�eՇI�Ĺ'��lN[?.-��y��x��{��E?U��]B~E�\�j�~����ȟ��2o9�k��\O��{%*6�A�/`�.O��l�V�LwVa�刅BB@�k�1N\*���� m����c���%�U��(�2��
�C;_�s��Y&5)���O'w��7��H>"�[+��Vĥ�e���-+��@�UV�[x�y�%�VZ�6O��:�_�nv�}�������	�+_ ��3�e���b�.��h�W�3GR?h!cWn�,�P1i�i�C����*�w��ۈ�]o�|��K.�b5��+ ���[�Y:\D�Z���rl*Mi��K�S�muH�*8�^L��[{�z��Y�Ap���N1�0�Lr?��	�R�^=w���Ʋ+�I�uk�	�WS���Cɻlc��(� ��|��R������2���l6�@��0��G���ޔ���w ��(�=�1�q���A���{�X�y�R�M�Ӝ��U�r��8��t/:0� �Ժ?�C�}k~ܶW�Ì����H�o��ɨ5%����X]NQ^@���z䟷��������=/qm�����j�A��P�]G('�����7W-����X��eN���f�"��^��Y�q�K��t���Et��˕;�0�/�ZLh1/A��;b��F%�
K�˅[�Լeɛ����jWŜڔ���Cy�`�=���O̦X*��#c��H��c ���CƧm3ox��#���N샽�(���%~���pc�g�.��/�e+�y�;�8K�� ��N��դ��Py��[�kw;�%���Ą�
^�.E���[4_�@�B=�eވ��Js�����ܦKJ�	ӘQ��H�vU���ҤZ�k��g�C#W$�ׂ�K˶�cHy$�d] +>��`��+(�����_�*�
ԏQ$A-����b�cσc:�xZ�:����:��_�<�/�.�Sf1��g:��z!dƷ�9t�ڑ��.��Q��J�]fp���+��F�=�w��Nf�c,�4Ļ|W��j�a����W�:�@	��eV$;�k�D�B��n������>��fa��o&��+�����/^�c��Ͳ���/���쿹!o��ZN?q��VA*�h�i��L�'���k�f7�W������������m����<�S�7i���;�È1��rw��8}1��=j:͇�5�*��E70���!��⤒�B|l�Q�ԛt0p� �BqA����j�N׆y)�����J)_UE��on�k�?�s�'�
�1γH����8��h=	��ªӬ!��%4lG��=�U�c۷�{}�Vv nr��{8ܺ@eet��k����]4����b�I��"iVe�y̶�a��S~�V��r�}��t�:� ��� �^y0�=K��6�#k 0O��eX��3B\�gxJ�|.+�5��,�v�p��Q��]tJ��A�؋�d�2)	Lj��8�G;|�z8����9&_����&�v�SC�ā
$����o��@4�]�X_ZX �i�}��PU>ta4�c}�}�'o�e��ͥ �.D{�Ԕ��OҬ���`-���x_���q��ʠ�U��t�}��vwH��>2��4������m��v�ݍԎ�`"�R��O&GO:Y@��!tw�	��$�z(\��S���E��x9���ML��*�,�1�sr��\�b� ��� ���Y��1~ynjb[YUw���:��Iu*(��>Ud�y�٥������*�W�aQ�u/�*`���#P򕍂d�۟�W�����>��@;Lu����gT�^�x�p-~���S[0�@h�]K	+B�u�	�i�pS�?^8��*��A�k�&!��Ӽ)<*�	�No��"[���n�u�!��nWI�!��zA�D"i�~�<̼�۫�)�&$����/5�^{�H^o$�H$�o3 �#���Ӊe>,pS�G��Ώ��6h$>gA$��h��:e�,-�R)��*	VElSR�������6I��B���h�`IsJ��B0�ˏƑ.�|x^�䭼����24�������B+�Ƙ��o��I��^9uE�q��S�Oc��)_��H�:hFg��.���������o�O�U�s�a�#`�|�D0 }M�l�;,M�N���\�X31�K`�)�r�N���_%���@(��>�^�A��,�_I2��qdƢ3$k�w�(�kl�_����BV���\'���g�i�b~tʐA���1Ʃ=���#��'��TE(�#��o���P��/:c�L������{����ؓ2j}�A���o�U�����9�9��AT�o��s֋�����$�w�m�|/	�~�����Բ��(O��:��
#t�%���%�fG�b�kxK�5#�c?�YT����
.�C2��S#ö�}�-���s���2��/h/.r�&w�tumEޞ�+g �Q��p��4�k��m?2Յa8�D�Q��H����\�C$��!;m�>�Z�2#�%A!T��T�o������k��_�����^Tk
��X0D���EØ�M��QmH�6�5��a�{��p�z���)�v�O����\������욦�3�D���$��r��Sb�9�Z���G^���nS�\��L���V{RN�3�P�x6C<�?Jau�5�E�5o6��2��
{�Ô#��W�+�WL��G��a�v!z�	��.�`��܄\bس�ڂ"HV�1�U��
pϭ���܅ѷ3���C;�ȏa��XE��]������a��Q��&��7�:����ZHղ�y��.]x���1�Md	1aK���D��Ī��fN��'L�>�D���
>��4*T��wќ������!�d�kP�B&.G~�f�}m��)�R!K�n[c��K憯b�W���3e�r ��|y8�";Mؼ��~�Cn��������ò��^��"`VY�\���i;�Q�fS�i���@�dv$Ne%�;ݨ���Z/��+η��u�,S�t;��ϟ��xj�f��D���
ް��_�߁����>U��1�$dו3�����mK�X�:c�B� ��
|5����\&��c���#�|Z��ſ�����ŋ�oAԾ��D�k(z�ѩj8���25�E%�����7q��������Y֭!�Am��o��a�4�`���-N�䟢��v��U�-���6N���SU���>|���G�6\8/��^����'yeC�瘭+R'	�'�E3�ҍ�����w:LB��-)3�>�	��kz������˹P�I@�b2�O���8n����M ������K~��LCRidG��>�A�lx.z�Q�?�ay��P���9Ly@R��O����V;`v��iɣ��%�$+s������M�]uU�f�J_u�"Dݕ���1Q��D���{u7R�4S%����b��F���c§�x��$tsJOvѰ@!+��.�WXa���b`E�z�Û���\g<���L5��
�4�a�*��%���eę�!��<��I!k�V>N��j�T�x�����a�z�����fy%�𫔿���$]��f/�IH�!����׆���Mg�����RMA~#ݞYP�a�O{��J�d�t~cSsX���;=���[�%���/D�?���6��Q#Q���
v�AuY*�@:5/�c�_wP�����^��(��o\[a�L(�Q��n,QȄ�|���8�xOq��oR�u[0&�<��6:�m�d���	���7� Je��	�ˀ��ɇ'u��>�-��S��#�̱�����E���x�������Ք>E����k�S1'��|���E��(��sx�}���TT�'�z��>U��ݩ�Fј/���b�0�PҴ������n|/kfJ�Q�!/��;���w `/ڰּų}Lߟ��
�>=����r;ț�||)eв�M�{n��d�,��䫞j�"�������P٭�~�	/HX5������3k4���6 �ֈ)>�`+szD�f�]+���;Q��ܬ7ނr��A:���r��;֌s⚏O����cirH�B՝0>!G�O)���
2��ѮnlB<%�E��R*V�+�W���Vܥ�#��ӐM��k���*)�,���x��:�,e�+�,�r�� (�8��]:��&u��6R�#N�� ���?�-��.�e��Q�E��g
l��Le���q܉�J�B=��Ŏ: �yc���<���:�����ZA��ڑ � ��cP����j���_/&[��8�0�W����fd���iI�E�B�]AN���ܿJ�t	���Ի�`�� s�|�@O)�&uf-���FA��2�gco�iQ΂��\n��D<O�S@��e�"�k��z�����$�tJ�2Ę-v�<�� H��Q�g��:.���U�Q��P����}TmҊ�b�+�I�<tJE�'��L��������\3��c��Θ�p&�1:rΎQ��8յnJ�%Q����(�.'�e�hB�����~�f��3���ZX�����u?��d��ɱiPP�C��X�tM3�H}��ć�W�	��<�j��S؎�	C��;��3���1:�ix��V�P��G(H%Ӌ�T��`���U�9�vJ�(V)����k���1������7�a�k����U��q��b��W�����*7�\ 3������$4�5;�FҼ�#�k�RdɂBl��'BD�ўq��_��¤֕��*�r�~�qF6����}BlӐ����D�`5nr3�Ս�Q�H��؄��s�%̛��M����U�F�;��:+��%�U�
���TomAR��\΃�W��Qi?�C.�|=Q�@�B�#	�����V��>�U�_B)Y���Kc�K��Cx��~���18S���O�w�
����A6�8rYxy���磜2yH~�z	,��BN�X��}��V�:?J`����0���+������'�2���g�u�j�k����U@2U�ѭ��Z{�����l��X.��&�g�^�{��92n�ֺ�����@�n�R&�|�D_�'�*���k� Wn0��d�TY� ��İDZ��rE)�<��9�̅^����!h��/�@X��G��ʜ���JP���8�̺�6�u�`0sp��o㱫��چS�����.懷�	�h?��*O����P��ۇףYZO�iK��ޟ/zcX�y,�*�	�B,a9�j�,�;�Sw%�o�����o����xa|���b��i�b��^RP.���[��$>Hő#*e:��Rf�=~��Uv]�W���E����۩?��:��Lc;A���a����cL;"	��F�$��}��[ !3�`�X�P�M��z��Q^S|�Q����%h�Eڗʿ��i3��w��8ɭ��G��p�	�z
�O!�ּb�������47�R��3�ʮ�C�Ny�X��9n�
o�s��}�X� >�A�V)(�L��ݵ�ĩ�|�S�?5����L >*5u�&�/�ڤr9r�0=�$)��Ũ��u��i��hl����R�.�f��ۜ�W]�V�f�R�>Az��3�$���?;;��)M��t�!f����q�?4THw7���������,M0�IS�XQ:h�hT�/�rk�
�p��|V���J��W��E`���`pV�m�Ĝ����rp0��c����ug�<0X�Dz��ջ��v+!�sJ�`-4Ơ�w��p�
�J����q#i�?��av�|1�����X�Q]��Om	P������I���K�֚7e:���44B��3�L�y���h<&�jj�un<��E��1_��_W1�܄|�:�e��x;ƉM*�v;�*
���c�Y P���q�	��{��6�ESM���Q���m^a,���]`J���9�m� �5�����{D�g;b�cUM��4[*R����]�����%S�[7(|R���gl�
3Xlg���)�p��:�
�cB^�t��9���u��y��t��:"����'�T�����m?����[��LPS�/+�o�m=�,H��k/]�zW=��6O_��
��}f����\�cC�2���}X�W�&]�]��Y�ώH훺H�S\1��=X�̎�ҊM����ʸ�a]���}¶H)���m�HDh��N�=4/y���c�'s�e����D��9�v4ܸ3��}U�X�i��{M��k��j�V��zN&kx/Kc��0��M��M���}�Y��Qsۂd���p"�Zw�Up�����!,�]�V�E8&"+ut�ћ��D���޸�e��)~��	R����+o7"�r�������"x��%a��P2����pu9�N��(���Pw��&����wM�O%zͱ�i�b�E��0U��8��0��_~�:}7.Q��S�s��j�j*�O��7�&���M�����O���К�P�mpJl$x�A�&h�QЍH�*i�Ny~�*Y�F�X����uw�����d���o{�c`"W����>�)#�6���^���O���Ts
�}�o0��%FF������}�ҡ&��o���*�tg,��XW ��^��|�D�tZ��-Bh�Xѻ��1K��j��gUt�k8�?�B�Y4r�v���W �oL�� �v7�j`Afh�7�j
�E���E=�=�B��4F�kt�	�(��!8f|���O�>K�����%�]7y������:ɗt���IΜ=�%�ơ^qw/�?t�P+�@n�+��KjN���5Ki��5���T��6"A��Z�L-�<�/tʰE�[z Y���1H�'0�;p8�P�U��DI�tPy�f�#�g�J��X���L%)� �VI�p;d��bu��[��)*AZx]�����DBSQ�W]�L
�N��n���L���5a��&�e��.#~B�,�Y��nij�u�(�㏰F��8��S+�y2g��*���B3�gW��N�`fS�V*ㆣ�z�"E��c+KE��1Ãt��(k�_�ZQVj�x�٤�p��S%�	J��j���I�sJ ���*��e���$[��?�:D[��5��WTy�~hП-�@v�K0��4�-qd��i����Q�yAE/1�<�*l��?~�^�/5�$�S!�i�(�G���\��y#��% �����P��D�����2̅	I�Ov49X���@�B���ܸ�]�/�=���sͱ��w�T�/�ޮ���k�Z�4pJ-�b�R�wXX-P�tH���e�b�A[W$��e��ߌ�*�
~P?��0(�n�ǜ��ujT��tU�"�h67�}Z;ZP%oT�w�$L}�ߑ�S�j� ����o�\�D�p�mx��X��u��
�z�6������)#^�LBϫ�Z��L8����f'�*2M�3c9�$^��D���鬓��Q.��B_Vh ������\��`on�N8��Q=0Ѿ[�W�����^3i`�/\���,�~Cɸ��2�Wx*ט=n�n�A!�r��WK9�
�ۡ���mY����)}�@</�M,���$�_T7�l<����&�0�P`���o$��G�ٶ��?�3�)����Ke�<�F��1�t\�ԮT&�t�Q�WD�����i�w����w�d	���[
���:C�y�p5�CD�^w��Tj������G�g��9,�<��}���tB��SWݒS# j�+"�7j�z^�u�k��ȼ\`�bQ��b5�1|H�+�8�
���޳����S��uO�6do�G���s��/��s���QR e�0��s+���𲨚��m���&aP��F�!t��A�;���:�OM�����m��|̀�wR����Y���q!?l����w�ֱ��� �2L���H&�rAf�O�E�j��qx���Mo/Z�_}�ؼү�Qǰ\C<�.�IuT�ss�v]'�Hk��XT�O/��(��Vb ���̈Z�~4�0�K����� ����ǡ;�[�ǣ�ۍ
�/����xei8�ּ#�*tU@"S$���F�J����+#\���U�Z�,�7�UF�&Ln{y�D0��k �my�q4 I�4���=��P�pk��c�e��Y�Sχ�����:�崉�7�?�J.x�
dz�K1���֧rC�q�1ʭ�D���:�8z"�[q�T��[?��ٌ�����˲h���s\s�O�8�Rs8��7[ΐ	HZ����[����.U�3�eo�2���]�B�+�EA�-��h'߰؝��9i��[>kT_Yx`��ѻY�����S������M��f�$0�8s���,�Y�l������-�z3��q'�\�1�`�l���w������5���_!��w�I��]��/I`�S���q�>`2&G�A��%�!ه3��TS5f��l�h�SX)�J,��H~�_~���ι��C�ށ�P-�<�͵~���P3�'u��<��4�j�1�&����B�}��P��?�]��%�R����j�2U���Z��8|�����	�L.W�?��'#�!7S|7'*�*��G���G���7����� l!d�@,āP���D�(��o�(��T-��Ol�Ѻ}�'Za��T���a��P����}�F<��9�k+����q�8Bhl�6a�� ������l�%`��8��n��j-��w�M�v@�w82��b����G��M��'k����
��: ���f4�a�[�0�N�E����I�x-�6���<�t������6F�p��u�:�����5S��ʧ�M�-P1 >8�>$$��F"4UJ��{"k�	E��s���r�G5f�2 <�� Cܩ%m^&��O����?L��-;[5#�}Z�܄f�j<|�:ʲ(��nR0��gu�A2�ц���N������8�rBO�P�!XY���uǼ!��!j�W@�II��޲A[F��p���#e�J�c��,��D���]܊����5��䅛}�	�~ �Ц}V����g���4gb��W��O���ET�]nwB�<n�sX���+���S��9��:�l�9�n��,�������t"� Y�*(rZ=��\�����V��s
�G��7fH��R��2M0zT�1q)�����]EH�h6p��ǂ���5;�� &|��ˏ1M�EXIj:GT�7x�K_*՝�l�!D/��B�y�B�G�R9��?�'���rV�Ռ2M��k��Ը_�X{�וhX�o���xWLVó;̯@y�] ���C�qᡓ���-:��L1Y_���z�')[�;iKm}B��l+������P>@�����3�W�%����['���<`)�l0�Q?0�SL���sE#����F;d����C�C�ʄ�cE[>�e���/����p��;���_6L��ڰ��_>Ǹ�3������lc����z��P�� ��� �\�����L'YǤY?c���d:N�H�z��A'ckd|[��#{�J�&�\��J�Q��f<�x�,����%s��R��8&��{���X���l��d:�c��l�Tl06N_��z�D{� �%&�Ңzm�*�a�8e�9�Ӷj�l��(Q�5)W�$lK�����A���C��N�����ʘ��M�)�/u�@��/��s��>48&gr�{#񟨸���X>:K̘0������X\?�g�Yd\ww���F�y�=���c}s���3&�c �$�p��\
�&�٘*ש�᧱���!^zC�4T:NR]� �����E�(o��!F�_�E&~���Q�)+������b����Ly�IЩ�
e�"��z1Tr�l\7iʆ�KE<�IG��� ]�m$��^��׍ŸGFS�j}-�
"����M��,�s�T���������ݠ�զ��R�^�����d)��<,�L��$1�'�h�J���>�`i�27@��#�<�i�kG0S�Q�m�����b�-�w!����{���M�U�^�E�_�Ė,�����.�ݪ�$�����Ҳ�yr�V�[e^�c��l���J2�@�u�L�q�a�r�\z2�ڂw��]���%��6rm|���#X�t����=�RH���7���u���,�D�%ѡtw��sz�ł��հ���X�pRo:T�s1��@R�ů;����Rri�o��(5TK��¤�0�B���qˬ���P�c�Y��o7�~�[�6K�t��^C�������{�;��}8"nw�|��X@�!��$,Oz ,�a�M=���f�w-���-Ĳ=��[����k�p�ܳP���-���}0,������Iy�@DjJTh{�ǰ�P�GpY	�$��)�_�>Q >�����@��T�q>HW�b��Ɉ��rw�𲥊��%�I����J(�K�n�ሐ1�|j�zx�+�c�N
-v�����-�\J:�9!X��-�����i)˰�`M�;�+��R`IS�A�["�9�W4�H�_���jF�!E褪���
#n� ��V
Z�S��ũP3���t.ql���B�F��<�Ji���'�HZ��H7����՘�
SgP,-�����^��Nw���|�I!	.���0�W�9����I���ku}]��e�'6�i�׀0?�u��+���8ص��DƋ�Y�����c_ѧ�?�֎[�v��l���*����u'	:?Ƶ)�KC�߲��.f��Z �s�vȯ7ςZ���D�������bKfڼ�Hy�,7��|+7��/�r��x&�Twn�x���r�]�;�����&Τ�l���(�rjV:� PI�T��ѹ�8�U�Dnէ���Lb�"��!S���$�Sk�K1u��Ō�\��i!���J1�����N�g�����1	��X���$T�}X lH�I�3U}�^��~9?¢�m;=��#���$�Ѫ�!�#��G���In�j�W;�ڟ���c�z~�绩sV3�5��D��x�{��;�C�	/����x	�	��X�JOx�ӁhO!��Z"8k�_�?�O22w.��14M�r��&�tڜ�Qk�ٰ����ɧ\�
�N�����q ӎ	��
���5�89.����2-�հ�vk�&����CIkl|�M�W�+��͘j	u��=��(��;8S�m(�9e�1�۪۱�� ��)�Y͗��I���)	&I���\�D�ȩo�[�p�����p�׍�����w����{�J�@�DD�ϙ���~c�O0!�\�3�P9�ўr�Zk�1�3	�秳�ݼ!�#d9a���h���	��b�\����kw�0~���7���C�}/⸃S9q����
t��.aq�&�%k2��Ȗ�t�K��h��� ��>ڋ?I�l�p-�  (�qG�n
ʵi�mһ,���N�u�`6\ct@�чA�ּ&�q'�FEv��)�ü�	I����'d�9..4Ni���"�"��E���J��
<z��v��^6L�4� %> ��z2�'���B��,��~�#�J-��(6�,�I��EY]����52�0rmثx�s��4����v�
���Ή���Vxt\D��ha	���I�Z����?~,���?�0r*V��.�{+M�y�v��HM�`<Sp�{�+��i<
��.*���B>+�|��M�D�y��MU#>�;�Qm.�N���~�����zg�r]�E�kX�>��Z*�+���^W�3lH: g��l�Fɘ ����MY,U�'Q���7s�`0�IgK��E�$l3@��[��?�\-�dc:Qk's&�nW���G��S,>����~1��8�Z)Ô��.��݄b���6�߻1[��!/��Ž� ���8�00�v$䞮8Eh8R(��|ec]��(��!d �S���|!��������}+1
 ��?���a��'��ry1Rrwo��]T*k1��H���-c�����P9!М�Εo,�V��1i�kR#b�D�b�T�L�00�GM�G�Z.��	��wK�@��̸������O�4J���R��+Jb�Lۧ6��|+���7�K�.D��V�#]1N�\�Ȕ�� ��I�\�{�ȜQ���������=5�9����8�i�I�<c�3�7�hd3���M�h���(>�?���[g���|���"^��V𶮡���L�!G�Irh�(���1I"!��DlM���&B{9I�,�ö���iw��x3F���%�_�f�%K8��-)w�����YY�%~���m������j5Ud	4Հ4G����SY�C���wD�]'�(���ŷ?�8F;�r�/eG��<b�~��kto#gl����cw�-��(�a߹?��۲�m~�6ۧ�T*�xi��0{>$r�&�4w����s�\�[�k�6w_5y�`�"*l�*�?�C�z�Ͷ���ɋ�\$/�r��O�5�+K��;@]�󻎣:�$�3׎�4��v�H@em��	J'K�_���kQ�+�p ��OB�����hꍤ�U�`��u�)pya�Y�?�\bJ���M��x�KE�Z���G(��*rkxB2db�E
L,j�$�Y�1*$&{Y���m�<)��|�Dַi���C�`\�/*7��1�h~�%AM���щh�J�m��kˡ�W��M����ykH��Qq�
��-�ذʠ)_��^���g1{O��0�wµw0���]E�YH�D�K�V>y�������14������͙�Qt����#:�r��ڄ�M5���� x9F:�9P��y#���+r��LJ��G���;X�{��.�����d�9m�9@CX,��T3xg�W��D�"?�L��.5��#<���s���X�ʊ��VzI�m"���0�/E$}2e�o��*4�CM�$��ɹ#�w�IHա�X���p���:B�}/ϯ&C�no�uE'����:�]Z�>N�(�_MZ+l�v��s��>�N\1Yb\�$})��P�poԆ9^'��Yt�"��o\�h��D.�աd �%	B=��D;i���c '|!�^U39	~7�x���kK��B�Uȴ܅_@BE~O���L"�ab�I�`�`T7ZC:כ��y"'�tE�TGu�Hqϛ����	����M�e��{�v�����tnOkC�G%n%aR��ˆ0���I�/1:��/�#��8qa5��3���F�w���<�x=w�Q@5_�������@��fy��n�Q�D�	��K-�l��M˕`n�7�È��29�0�����q��!�x��>�v��uM(��2E4{J�{J�����B���B)����A�A�º�u"�5�
b��̫�(���ԩW��fz� U8���[	�[aT��AA*jK���D>�	��>H+/�a�B�<�(��^��1>�垖�1�qU��}~���~������rw\��/���M��#;��K1JD��WƊ�w*�W�V���O��t$w'��y��)�o�D5Tݖ�0��X!���<?1IW_~�W�ܟ@w�o�g�<��T#���(�Cj�Th�53S}����gw����P�8)�򑻊X!�7��%R�_�g������n���V}-�VKWj�z�
q+���B�� "����*7�����3/���H�U������Q%L[��p|�QHY�FЃ)ϡ��>�Ԩ1�M��8>�'�-���e#܀�!q�=����^��fBpP�Co�_�J��Sc���bC�q��[�z���f���P��-�� 8�|Z$G1�O,��^Q��5#�[�!��XI�?Ӂv�|�[Q����5��[_�R)ȓ8=�%� ������O`�St�c�y���b�w��I(U,ڞ>Mj��#g⦺�����f�¿���(c�����&�Z�r��簋{�O�����WY5�W3��UwP���mB� -���k��r�5<[(��訠#
�4>�9o&���x�V-�bb4��$i�Q+�Y�;[�&�2%{����4z���4�XM]����^�XB�W7Jg�?u�y�L�ȷ���X�|ʺ��Nm:!���	�ZbpPz�nO/��m�k-�.� �p��rw&�'���*��r��<|�/����/���#zI�AnU��Ip>G���a�Г|*(�hc���`�4@p{H�6M�D������<Oer/pN��m�]VȢ�bN��y�n��i�*���䵝\�0�u�7��|����
Β�z=</@=$,�L`9���1���f�C���C9���S-Cv�R���������	�c�%�n�Q*�E;�l��w�/��#k�u0��Gy�&L�.-���{vc-�L����b+��.��M��MR��}��iMob0�5j�j?o�V�X�������t�ⳋ
7����t� NNt�%�E�bƴq��+��!L/`�:���x��'��,����zd5��2��~'uС���Ak�Q����{UIABcw�0S���4E!&A#��>�˾�׮��3�F�U_+�Œ�q�����r:��ӽ,�r֢��d�5�Ar�����P#�3�|?�k#l�Ax�D`��L��6�7���^�\^�fW��&"PA_-=�����KDA�	��	N�&x����UٴS�)�}�L�W��Oݯ��g�)
��3Ul��c�Q�Z󵫝�i-�5OiV�2+*Į.M%�W�#��*U,��D��Tn)�:a��$m@3�;F���ZF��?g6��d�W)U�;R�d�릶�a+d�Tys8��vV��n���|I߄�T�ڥ�9�,G�ht:�W���
H�)4�Ȕ2�ƺE�!7V|IN@�iql�PPځ�Mdu�|�o�,u��Lޅ�Ǡ�@��i��&���-�8��5$-rTܷ R��W��c��q'�d�����������?y�ۣ��3�f��+Ϗ�6���}�l:g�4H�-�f_��ʄ�q�a!*�LC.�Ӌ)��ײ#[��|�����+���_A��A�Qz�����P�Oj;!�nOZ��I �6������(�i�.��Q�f��e�վ����FV_���R�;����AW!�:zuH��)춡��u<��ۃ�E�dA�lQ������,nFC�n�/���	w����o�[<ځd���RZl����Jg%q�kOX�B�x��Qtcl� �s"��
�R��
�@V������A����Q4�j�t�ʦ�r����,RyѼ�,�i���X���=��mCB���[e�i���ɷ�:&�b	/�Lrk85I�Q��^�a�µ�q��q?��/�����\F�̲���/�Tifp2���$7���dԜH/�Y*���WB�kh�� ���X�B:�� �j("�h]�:q����]��4'��I_ܦ]F�jۃ��sG�Lu�p(���ꆲ��}�U��f8Ꮶ��b�����B;i����������������Z^I� }���T�ǽ���P�1n;�p�{�S��9�y�fú���>NY�jM��b�;�ĴZ�_�MN����^Rrr�����WH�	���1��o� �r���g�ed�I��� D���DE�H�2w�̪��,\"�g��/�ܡ�z� ��i��T�Qh�����s���>�RX'�Oj_i�X^u����#��Pa�.�{�|��]� ��� ���U�5��Z)�GZ���9y��oT6�x���L�Q�q��I
�اM�<9H�!��"�3F���Hw��xP�H�n��V�R���۬�$���q��돖��
`i����[�q�f�Ԏ��(ݪ�k-zXt^��tE�!�KL�Ęq��#��u�����k3���ZqJ�ӿ�I
6<���&���o�������jn'xE�Z�av����Qx�gmYzvxFl���%��̑W�#8)	�r�JO�Z����(5�ӝ��=�������3��[��ܪ�� �>���<�C���Yޭ?!X�̯r?�����d�^�T/��#T[�3\(*b��J�,mAl\��R���{9��[4�-�]�=�luq;>�����Db��bA-�ߪ���?SH���"�i�d˄�1�r�l�~�O>�wu��5X�6�p��G$����l��m���M9�^�,k�g>�����_D���B�SL�.��[��b=�Q��D�FT��~h�.�?�F�i)�ޑK��u.�r�JW����Р̍�e���}��_C.�+P�jx�~Gm� �� �� ���P�G8БN�UcվYU߉��K���&Z2ˋ��2�=���gy�L�������G��z���A���=/͉$��̾@��h~J��HZ�R4�`׋���X/��E����4��+\Z(��rV^fd��h���Ix�t�Zߡ�+2YÍ^)wx�<xZ��J��JV@�;]A�a�߶Ǝ�Z�A�7�D�u�c���D���!���Z8Q�l��n��!�D(��*��Yn�$�}vW��ӡ��rM��؂��-Zf��M���o#ID|��ߧ%9�1�}��P6ŷ)b"o�qr+��BHM%2D�^�;�G��Td�t%p�+���#�Ƹ��Ѻ���8{Yy����R��bm���A����\-y��C&-t�˘���e�ƚz���m*���a��6��i�������h�ڈ��diA��+Я�i^���9!p������0N�vX���3�0�e��=Y	� ���2��&@[v�h+-p�0�Kϝ}�fgZ�0�?-)A&O�*V	Q2����Ч�4����n����si� 9�8���84�=uLaѥ��e�)J��-"|�e�p�j��K�|��z ��z��aPY��k�`���u��tH?7�#�ix�S~��zs�U�_
�.�dh+�<���cp����x���]��8׳x	�����Ej˽��g�;�dV;������^��:��CH�]@1_:�o�_�+��#�����e��v�g�k�V�!��=*=���y�����6~@��O��]�|F�!Daa��2A���:{����>�2x���W�g�Kl�W%�M�b��Y��nx�T�j����!s���'��04��%�KӃ�\�O����L���@���r����͑��tٝ3d,QM۵0�8uWI#r��m2���̮o�m��A&H��B�&����X��f�+*�5��q�s���(PV�μ�Wq,AO��\LAo�}������Jn�sH���?k�;��(���y>��U�>��h����5� 
P�����-�;tr9raE����/�tc�K���x8ǹ�&������p�ɉ{툼������<X�g����RAͳ梵=5�T9u݁t�s1},�=f+���6�$hVm�f�����=p*�����=d�ڪ���n6���굸$�\K*��]x��ѵ��B����6�u� �y�8��P3�CAgɌj�Q�7ғ�O������>؈D6[��@�O߁�&	x9�K�w�a���C�|��[�|&>D��}J�Dw>vj�;��ֻʆ	U��^���铎�%x�����"֣+�l������iK�MQ��(�w���k|�|t&h�E�]5-�-��ɶL�v��ikwJ��<���[�������L�u}�)�b�����L�E�«'t~/֧�8$�S�4����0 Xi�`U���y/���7�Ȃl�z��Բ���<�(���EL�#�x~�~xK}�Sf`��r(*�^�����k�o�L��N+�����v�[��U=A��kLC ���u��]�K�tho���V�5��B��ֶ��~/>��t���g���^.��Ѳ����s�]�|���^3ut���=�ZL.5���I�������[��E\�]/�^��m�aBnU���e�dgm�ǝx�)���-�����v�e>��F�x�&!u�/C����W�*D�r]?���?ɳa��7���^��I�o���HCw�QB�������T�D>�`6p� ����K�ʰ��l�\N/��IV�e�4�?Lpc���y���;օ>e��8�5Q��4�3�A�X���T�T�
)G�B}�(P�*�ߏG�-Y�Ch�\c�
<T.c�Z�����ʕ���,������i�
�i��oYiwD�Gh�h0�2-�砂�滛.'S8�����4�*m?�5*��y6`���N�{�8� J�"�j��C��,��_��$%���}�P {��)R.�5��}���~�ST�4򇻨�KnZ��d/q1�;�b�恝_I����^$��[д���Y'���W�{G��e�D��m?���8��(=\L^f�v{D�ߍ��~����WP������_;��G��%a2�7����
V���������qh~d�����`{��L'9d6]U̩�k���o���o:e�C����Q��jkcR��VX��r[fsZꯎ_U	�`�V���t�b4}���7�)AQ��1��1���Ӊ5y��au�:^=���'�x��	��z�}�d&7�/s.Q�p��r��O���,��Q�փ��v���:��:�"e@�p���1M!��SQ���1G9��>GXf*������~-�|t%��w{������c��+�����E���.�B	����	�|�� ��`,��H��е��ыh"II#���˼fj3>�=��Ef�n�1Ѻ��ch�X�@4���:�Q�Z�S��qֲu_-���n�����k�o%ƞ�Q�F�-Y�/��q�t�#r�+�\���\�K�]�
��B�V��n�V�zR���a��l��ݞD\��k頌�%W&Jy$|:n�Jh����Ҹ'�ɣ�c&Q�������\�������=$��<�*f����<YV������<�\7EK(i��.R��?�y�ʄ�Pb���wQqp߻[���J�jtSS(���m�#��U)q2w�,�KtY��Ɵ�-�^O� ,ߖ���朗����N㬬$�r����E�I�r�C���'���0�O�6C��|%����_Qi�7��O��lZҙ�P���֚�&"��t�*�����}:�Z ��������|9���u�L}N[#�5�m�����:<����Tv����O@�}�r;������N��D��n5s>����eV:"���05L?u�����]�����W�T�=Jh�.K��z|���J���2����>u�0��2�;�Æ�We3��=��r�عԎ_�Җ��8sx@NxD^�@���bB椷&a�3{�j�eÎ�]8�{�Xqc����[)����G��ХO_'�	�`������BG7��^d���H�ʨ�LҀ����.��<)@F@
dew�CE�9ż6�5����`+�]���k����gvPoR��q�����s�#�P���qy��G�@ Ԗ.$_>W�,�q��I��0�6;'����[O<{'�yt�{8�7dcW��L��N��"���u���N��H�U�,u_�2�\C�ؗ{g�Elv.��$Yy)<����!����c/�x�Sy{�fYDSR��\ےq����$���%�)����;+��Ava�v��o��	����"󓖙�� ]I��S�N��ۡ8��$�_r��,K��M9�u��K곥� ����DV؈���*����E�:���vܣ&ug��L�;kVi.���N[~0�h��M1�Л�6�N�/�F�7�ȌJ%Wq�ߗ���/��?����Xt<���:"c�����QD$ϰ���L�j�fwh7^r����e��l!U
9�:��ۗ=9=��k(-�sA�3��-�T�ݿ�4m����F�{y��^6Nv0D:c��X����_�Z���[Q��E�M���!x��|�3J��ʀ&�5��	L6�Y\�#�6�/g�n�6�2����=����W��,N\�d�I�?_�E���5��6�����AS6R܃2*D�Q�Ҧl��4a�������8�&�-��w�r��H`�5=c������ƫvؼA�#���j��)����W�h`��ak��=�W����gGM1�����PB{�$!�mZ$򪡶����`��T��0+�#�O�7�ǭ�5U@��&dj�� z)�_]�B�^ĪJ��B(&y�l^����~:���ޡ���.�yz��<�+fk4�	).��Z(�iaPq0��j�y����'J�0K�����	�`9��P�GM�]��>a�w���f����$�^�4U��CC�Nч��'Γ�iA�߿�)=w-�pz���6WY5�}(*St��k��(��)�2�,��������E���"@ap�%���kV��"�o����&M��+W��/�3�h,�Oo,r�^�8����)AL��eۗ��Rk��|W���bO|��� n�����6����G�'o�1�zQ�2��k4�1d��Gq�6IA�[�ףȦoc��<fc8"��rl��#F2�
"��99z��u��je�h9pCs͈������b-x�3 ��/da����������9
	SZ�D0E��G�m��"�$����kG,A�S�GE��M�FY9�]�8b�����`mejC|wW(!�m�;{y"�"/5��_Ý5^q^�m��˽G�$/�k��/���p�C�ٮ9v286��P���U!`�]����g'���\ i��ө��偡�h�	q�O"Ђ�ܱ���h����ȯAb�{�&�8�VN��ц!�,��h���ΒF��Y�)a��g���X�)+W���8�x���ZA�G��Ҽ֏84r.Օɉ�������]{��	��Ъd�8��.ཷ�ǀ�%c�m�ti�^�&���%`�B��;��M@=w�ߏ��Au��m5a��pM��⭹v����ȿ��3��*J�UQ��4]��;]�y����� ڋ=�!xe6z���W����$�R��S=!��ɺSy*v��yH�T��|h�t>�Ic��U!�F��'�X�U�:��n�fLg�g��^�ϧ��|��C���z��k���3>.�2㚐�wg �WS$|e��[�ߥ�+��hk\[�.�F�%�Ҳ��6��&��~C.a�4qM��-ť�q?��~Z�T����!����B�Dݱ�gC7u&��Y�M��OLOnü�w��Z��� B����rS�B�.���`e�p����#�Q%�6�Eѷ��E#a��vT��V������+�,�����M�i�V����PG��1���Y!S���a�܈���f�*������� ���O!�^��
vǣ8=�V��z��V~ڸ�[��AʤwFS\����?Ѫ���v�'E\#�����:����t���F�Мuv(�ݱo��(�Jf/F��ۯ���l�ʱ� \GkfR���9��"�T�*��1G<����[����#V�ٕ�c���M���~�^޸"�)��OO��4��㿴{�v��eWUJ��;F{(�wp�f(��sK^4	$}K�D���ѽV@�p�|'�{�N[����-���~�:����	�=��^�V�S�b�0WRTh���d;����4�x!!@(��s�K����ʱD�	���B����7:m�e1Yy���Pu�g5�7��2AWՎ�P�H�Mr�!SozQ���rGG��N�X�����l۹�֤��*p�$����O~;��(����Z��������H��s]�PghG�Yw����^nf��^��ջ~6.���A�Z�|�^9I�d�8�[0"y�H�t��.�5qAj���g��_�1%\���g��	��i�8���$9�i��ǝ)ӢH�?��b��1���d��g	��ZH����������~W���ͺ�j��<�k���B��Ȓ��s%�L0 �s����	�����_�@r�|������V��&H>��*"�D䮅�+���2aC]���0�=cU��:2�(.�<�!���T�����,��f2��ue��3��hm::�A�6x�
mV��0�h  ¯���������0�(��j$���DY�CpT���xA���A�&���i�N����`��bjb�e~v�X���qvuz+��T�r4��З-F�,�w9=j|L���MSD�E�N�����"E��ɻI�3��u����$��"�b<,���\��0T$���ȞKl��v�ʉ��q儝(%�����K�C
|e60�����!!555���~�h�3�I �-�9���GG�� ͳ�v|��Wȩ��X���h�}�� lf�]�k����E���пr�+DW�/W�;�GE��"�&� +�z��fi&)_-��Ey�����8D*>�RծS0u��VW�ms�hҎ�c����ɇ ���؈嫉&�ȼ	�-19Eo�ڦ�cW�EI�7���uP{�%��f~��U&��Ɔ>�"��r;��[Tf�(���#�m�(�.��l��Eq+��'rc�o\Xx\�(��(��A��7�-OR���<9�_ڪ�~�r�7�8}s[�/���=ɠ`%�@Q����V�S��ǁ��� �Vn"}�C�s�[�d]�-!�Ҡ������sM3��5Z/W5]���O����-	Y=(��0S@�?� $�j��^r!j�s� sXB45<a#a'8�t�̼X�}�$�t��-�{���7����	����� ���*&�z2����p� ���U���.�RK�Iω�9��|��p�K#^����R��]׀Z~ `>����!1e1`�ӈ6�xO�����c=�O��p�~��ȕuO�n�|�;`�V���y!ph�@2�+��o}��4����1أ�D\��c/���s�:�5}�RsB�!U���HB�8�}ũN�]���Gkf����e��o���C�� ��:AopI�ц��I�g��]�kb��`����D�@�fDGq��1pm$����ب��z+�hX	+��V���bM��:K^�L�PA�R�0�>�T�����Y�ࣥ�F�*Eߙ휟|�淀�p���	Ɇѫ��g�O#�O0�Q�_�.2�'T�A+��H�K��N���b�Tw,̆$�t���; #7YQ$9�9z�1�*@��l�n�"E�8G��_uw���y��R���+W���9��\\&b���>����[k�
�U�����*�(��k F��r�]�}�v2�7E�A`�>N�m)�%��]`]�t�40�g�K&�x�O����6��*�{���C�MdN FD���!�� �i����)�� n���}̯]7J�e����IsU��*�������kX�
��E>(q|^q�|Db��ǔ�cv���A�l��g��I��2�����}.�@���̢����p4 1�A-8��ˉ��ݻ��H7�_��=_k30�Ģ�N���������$^��F�4]���
a�K����f��ߧ�u��}Kׁd�VFK�f/AdN�Q��/[����I&�h �%R*����R.`H��C�o�8��0E�MW>��4�zB
����R��"����>�r��C��񏖕5�����E'n�����䚥���{N�c�&z�G��:Z":U����%�X��/q
q��*�气�9G^1�D�,e�\k�k��E�v�JU'7�Aijk��Ρp��%�x�vI��X�sp>Js�>Y�8G)-=��j!��B1�l��w���){h�S����H�iDZ�"|:[/�\�2�F�&˺��Cn`ϗ8�c'����Hr����D�H����q	���j�&�b�>�&����p�m��Pc�6q�j|���t�d�ȫ��Xa�j�U}e����5˛ -�L��ݖ$���?�g��NVV��`jlk@�	�t����ף�!|�B'̀�m�(ƅ����^����%:�\))���S��%<��Wk��B�6{��sŰ`��|��K��&�|��z�db{��Y(b�	��Q�<�^��)��Fp_6D߻EM�}��9^h����C	�&����m�?�|PM/ƚ��X�:��}�@�(�=��6N�ő�0�<o����c�߫cH_�y���o��fs�5�kO�$������Q�![}�2��K5��A��y#���9]Ey9�ha���㕦�$t�>`Ӈ�����0 @�V%���>3G�F��W�i�{���hۣx�O�r�{|¤Ȟ�gB�E%ޗ��χ3��9[H�ӿ\�=z��_��6ė�+E@A9%�½i:>X��,݆s�C)4�����_�ɂ��\�~RD�&��J�jm��V�;7�Z]��+Z� �P9z s�?Z)k��Ƿ�B���9.J���u������놀\)��"T-'��mUu=�n�?6��gu����!��;	Qr[\Yā��Y���R��2�����i�F�F�"n�]�'2�c�h������#���@1��h��>�VX(^�7pu����U0�_^4k�H�+���sFV�#ͤ��c�v�4��F�1���ȳc�H��&�\Qr�v>>��~����\p�� �@����1�k�+�Ǭ,��� <-�� 6��;�Wr�"B4�$��]#�1[0 ތK�i֊�V�a�jݑ�-��	��?�fp���Y�_!�nU�{Ψ�CJ�����Ǹ)d�[��]��<�����z�pԤ��d�����D��| �rМun[q�a���`[xJ��1T�	�rD���dmD6��r��)55�) lQ�qp�T 9y���p}��>B0�R�7Ny<�L�{:吃���*�J�:S��75k�R-40Ç�"���v�^����N���TvȻ�oP�R�^�(ܨ��mO�ر�puv'?n\Iٮܿ\.f��a�+�p�^�e���
�)�T���G�hƭr��ӷ>��� $���0:.�;Ω�u�_��;d��䭫.���J��4$rG}���D�}�)��7���}k��V5�v�,y7�>�ę/O#U�1���&�I:����n�)�5ی�,���z�<�%�KEht��r�)u$5J �:�g�UH�����盠��@H�ͳ���Ť��X"�*���:��a?bi���h#��Qɧ*���bO�g\���״����*Q°&���߽9��I?��J��=�����kڨ0�M��� ���pC�ǏN�/.{Q�˖%��J;����~5ۭV�Ѩ�������D^A���꒮�Y��$�n���3f������X��H��wVb�om��='پuށ
�܎+��ƿ��I���8eې������4j����nAҿw<�	r�9��w(���<�>��x���&��bp�q�������'&l%�D�F͉�/	�[�s���5z�*ZP��R���������2�}�F�&�x{b�ʛ�'Z�?����ĝܒL����s��pGe�B�A�K�!��*�O ��`�_ة��O�+a c�g+lY 4���[�/�U��p݆��&�4;R��|T8����yאds��)t������P�U�c3�v��_M����f�?�aP��`=
���(�k1}*Ԭg�����j0���<?@�+<��#¨`��϶�ҕ�ѫ�����)�� �d�&�T����څ����ƪzUh�7���@�BH|�sf%2qS4�~lw�$�\� ����W��{ګ\�˩���]KE{��;̊|K͏�������+1��1🟳e�ܫNs��g&�H�Y�5P��xf��W�]�^����R������=KD��tt��e~�>�iǞ�	�0�e��Ը��O�Zg��A=�P�ˑ������-H�����`%R \W1����^�4�µ�$�z��n[�ʬ`�(��h� �p���a�S����v�a�˓f,�J�W+!����eA(S�ޚ�eU�ܵ�%�a}v�k�FbrC:5j��"�?��p�鲽g�'�=�J�s��+�M����@B(/n��,&E�9��&q���\�����f�l�z���z��G"@���FG�M,儦y�Ȅ���t��1S��U!P�}@�꫋���p*f�pM�ʐ�Z	�п+p̻0n���X�X�Y-����������v��O!}�Z	Ky:�3p��㾌x�H�	.�"y��8TҞ�mxvX8X<�C��k����+O�����^��&�l.�����+6�;eӛx�|P�Xz���}3Tf�\)�eb�[�`ރ����d(bHd��켓A�]�FO�0��izJ��
�L@ag� ��`7�EnԸ�;FY����at����y�	0�B�T ڑ0w��vg����gk���U5��X �n~@]�����`?�4���Y�`�j�����B��ɭ���A�4�K	5Ǘ������m�.�yٱz��/֐�+���ॕ��)�zM`<v1��2��^������덦�.d��RS�bca#�J�����AE�"�r����S��S�ih����Ysϙ����C��մ8����Z�r�@ϐ��
�	;>�_��K�"f 5��k��CQd;�=��c��@���*Ē噱���-P��MR���}��ՀI�Z�P�I���3�:jK�c���!XO���:�Nm�>���8��a�c[�l�V�&g/�Aش���%ˣ��M
�ε�8�>���_��۴���� _�4��gTD���B��u*�d�B!
sIbΔ�C�p��4���E�����Rw���+��,�����6�# �O>��;���=j$#p(�:-{&,�&��ɒo��
x�n����}�mL4%�����e ���A����R1�-Z�H^����F��ӹ6/�a��v��I�2��%�����e�f�|�^�\`n��m����$KlCA^��&���tKOYK�.$����İ胫�e7���j�3X��
���\<����ЀLW����ǆ3����NA�. 5��Zy�3Ƶ���f�s�y�M�*G]�-Y4�����Aq�,N�����T2XI�� 0y���GD
9��U��m��_�HŚkY�����Z���R#-�ʝ�ȧOF�D"ǠyK�-6�L�:=�wqgA�p��	�|<k9$�Z�Ö���%�~Md�MN(w;Pl��
���K�R���*�x1%35�Ņ�{�=����k�qyL,^���FY}�6TU2S�|5޿��Զ�b�;�3��WF��ԉ�-��!	���4�:����:q�|�]�`��Sy�_�I���t�t*�u<_f"D��٨��r�h'�q��utu�6(K�!	�2Vi�$�I�B�� ��K��m�&K��Z�����k��:����4OD�,�Hg՗}��Z8��&� �ە�¹/��hU���Ӣ!�ω������t�w�Zs��b�4Ԣ+b��n(zh�H�.��TH�����ۤ������9 "�U.@l���K�6��r�,ѿ�2A>WXJF�H�)i(]�"�6������7���$����|gUQ�~hPwS�ؽ��M~+o����^����WrN4��3���S���{}:�יj-�:��Q���N$exX��S�l���?�!(� X��WCJ�}1���%UQ.}�e��1?Ku��vuJ�A:	��>��	},��ʜ�Q� �v�J[Z�(��D��,A#�������6���f;�Ͻ��&�?Q	�xa���-�Z�ѿx=))��b�_��hM\�{٠,���>��d��<3lGɪ�����1�����\5"�;���٫��H�=F����o]�4ZiDq.,�G�u�k5@�88,�����q��>��@�V���{�TS�EI��V�%�=�}��c`�I�?�C��&E�2�#�`*ܵR�t��TFH��R&AD��$�YAo�{��B�*�Mڔ�<�j��8�C~{23㾾 ��@� l}k�Ï�g�Kx�K�6s<�Q#����N�[Π��z��NY�FH�#�k�>�� ��So���#�a���m��ƻ�m��f�.�AJ����ʸ��~]����4tg=��e"j��6m���p����j_�I���{������mU*.�A���R�w��$p�O��og����9G~�"^U��מj���u����i��]�K��k�����1�,�p�f,�NP�\J���Mڿ�{ǝGY��AH��<�.�e��	�u~4��U¢�<[H{e��p�e����M�4p�$b���C�0�ϵ'[�M�d��d����Q۾�(�{	��McJ�qV���)��8�1]Ɯ J��4�g����w�9���� U��߸�B�k൒M�tLX�a�rXU��t����y�0��\�B�_A>�x$+uR���i`�H{�� ��E�֩�wQ�9P�8�a@��)ۿ�xf�7��]�[51V/����ٰ:Ōy0�BN��I܆��?
"2��pkC�E���Q\�g��Rd�pņW:�ڛ�>xFG�'�&sA�NQ�g՛�25!]u6�eQ����ψ �#A��u@b�oȋ5�o�QN�de��ic��(?n��rn��f��@̆��]���}�W{
b�=�Oz���,����'z0��<��w����
�v�/��3f���'�j$3�!��,X{�C�"������?li�.0�� ��5d�9@�>�i)T�j�u4�5G�;Ɏwװ�,u��ar�!�NBӿ�$L�K�\���V���N�"�<�@��h�4�i[-e��)�<�iG��������,T�6������2D?��B8�l)"n>[�A�(��"X��w_@�]�����]�H��ܼ�Mlb��C*E�.h�vG��?:�.�$���!��ۭ1���j~S�Ὂ0���־���4D�]�o�e,�g+�� m���`�g�M7ӻܑ����a����y�9朶��on��;D�'k�k+�J��l�j��� �U�fc	��k���鲳-jdiE\�`C����Q8;@J�>O+�*�Q�<�z8�OT��b�;���4����h�yfw�nJ��PeZ�v=�(�ZaQܫ����b��F�(���{�gW����H<�J2AO�6A*�����J�E{m5��p?ཌ�����@����uP0K��)(e-_�[�!�'Zd���1R���pt������������F�&0�d6�Q����ײ�6�F#0r�éW؉��Z���������]��C�[���ΉiH �0ڈ2�<\-�G��%^��N_�����:� �^��n����0�5V�ƾ]�$���K�����"��� a�ݨ*8r-�:MV�Ȍ�H�g��oG��0�A�Z(�\AY�r,D��F����9>ͤ� .��6��Ѝ�H[�G�O�\���Z�#Ǚ�h��t����A[M%��(~g�|A&�8��_[*��t#1��	z��(�=Жj��gr�x
�	ʺ��湅S�B{1>����V2cÎӞ��D��6�D�EFei�ڒ̟En���s˦×�lz�&K9�ޘ�!9$mI�#��5����Jۢӯ�,<d)��s���z�G�����Ǔ��n���p�zQ�}N}����4wm�O咒V��	�ҟ�Y��Q���m\*�:1���'����'վ'=˽{p7f���"�,&�p+8!����C��_�X��M��8��� %������HZ���y1?'�xO*�rɈH�a1�ޯd���漑R�w��@�	"|��Szek�J'f�vX�� �V�M)�k�hث���}�f�tt��&�m ly+��\2�=BS{?J�f�n5Sw�������~�NL�{2������	���nB�����<�%*���y���X��RF6��)ُ����Uá\Uf>xݯ/� ��� t��&�o��ߡj�8�����:�*��waT`�z?<2r�[87L2f 4�/���[?0%�N�7�ƿ!�j,�A��?��C��v�`֦��ߩ@��)��i�c��fZ� �r�!��}��˰�����+j�kcV#�l�-	�hXX�ߙ\Ͱ�����������3�G_"�\����Y�"�ot�rs�<�B�<��F�r�h��bd��WPa���S���Qy�C�>����0& ��M�-WWiX~`����"�]V���?j�H#��@�tl���U,��A�2�{� �wKp��p@U
��^1���M���0�q ��?����+��l����D����!ЦtY�C�G���A���#8 
<<F�W��M{;G_�����.�?X�g�Io�mq{�c�,#�kg�A^U^#�p���&Q8��)o�,1��дzS�|x�T�.�\Uj���&%� ^{^�W��t�`��Ď�N�[�/e�X�Z����e>פ�T�׹ޫY����3_�ݪA;�U���+�y��=삏�����PP6Q߭���N��W���2��0����YJD,1��÷�q��q���4gF`��6N{����c��n�W{�8�R	�z�it1U[�n��wo��{�1GP� b�+�
 �㉤�SўUK�p&��lѮ,���Û��m�r�c����D۩e³!��gl:���=/��z���m�����Sb������d՘�L�9!�8j�Oξ���k�u���yг�K�0�w��+Sy�R�<m@}L2�r����n��3�����~�5e�R�+6�:��a� B��� �55wIO�s[��d��.s���I?
���Rs�ߢ-����c/���PV[q<q���q��M�~c�*���D@���#S`����:��4��F�
Q+�̔ڊ�c8Qm�\�d2�Lǀ���U���(Lb �hv�|]�1�dDI�$��]~�T�_
l�ywZ%�h� ݴ���G}�7�^�S8Q_���D4<��}7�eK�AS�M[�O�Kd��GZ3�؊�v��}�
?+f6+˧Ra�=!�A=���-~;8tPI��[ػ��a�Hhp�x�<�0A~r��ȸ�
��'ǂ�'����ݩ�,Q�п!��d��8�0���#�����DHox�V�o*���J0���� nV�w�1h���Dh��)�:xCj�@�"a{:�\�xW&D�,#"�������~���oQܞ�������6�o���E�L�N,	�.4)�����j�$$��^p�H�Q*-�a��DJC#����
�b�CP��Ya_w�ӌ�!�!�� ]s�EF(��	���"��ivT��@xW��aPJ�D x >�!LCG̏���Z�p��1�E��UHY��Je�^W����}w��8BC6����z;���Hr5�?E�d�*��'�)'o���\G�Oן����8�D��@<�[C߿4R&�d�2{ហw��x��b����A&�d	�\�rS���X�<���"��bL;��
��� h�K��T�L���9��R҄',�jխK$-KD:����1ؾoHB��� �l������C2�㢿{�Rү9<�~��!����P�$s�f��r�yfX2���b����̦�k�����Q�ȗ�JJ�x��`�
�_;M�>��!��u�85�AY���;�G]'H ��c���aw〱����9���t��D�oԚ)}J�����='6^���Kt<���8�b0��V'rf3,��W��E�n�B~�pg�ǴMp �w���C�?�}N�?�e����;����g��
�j���~�!Qu7/���ϳ�z%�R��u�W+&Q�j#0�����{=�SՕ�5}Y�l��Oy��	���r�T�pD��=��ڸ@�Z~���`��[`|0?�쬤�b�#��5"�`5L1��1TSeU�6����p�����S��6(�R�H�~�Mxy�����(��mq(^����4:�nWj)�XY�'�cjC{���8Ra�$aP��^p��F4�zp����U���k�Lqѣ�ݯ����$����y4&�L�z�a���~(�ȟ�g�'=j�v,���YT��ㅕ����8����g�}����&tМ��X|���mQjhORjx��q�EPm�v�̨(�/�G)��v�6��o�~?*����2���u��uk� f���p��k�I�\���f�u�
�P���*���,�K/Hk֩w Pe��y��7u�P)�I�\��6�x`���=�O��?�+T�U{/X��r4bVݦq��Jk�y#c��Fhzařu��Y�+�fe!��is�U���?�E&�f��}^��u�_�z�������6���
���MK|<�%ʄ�X;E�O�����Pˌ�M=�L���1���%B����1�r7m�eE��]�>q*���?
rÔ#��q�q�߶w�zt��n��=��&�m�����}a��n����a��iI���s����O'�_�i� �x�Vu��_\ Y�Mk����i;��m���t�34��G޳KG3�~�}ެ��]U�P:?�Bn'��#��#�9���i��d������]�]5(��)P� �"��;l7�Fn��C��(*傎�\�I����CO���[䇅+�[��h�yά���
%>�l�5yF�,#��=dd�g�L��q�˟�f�Z	�ކ�37/�:�'�KA�eT�g?�J�H��E��d�!%ނ�#8	C�`�'���C�uq���-��O�R��ԂiZ��6��}\�?L�.v-��Wӛ�l(F��ӻ�@�����S�w�X��7'�dh�?Q��'%F��#���4���D�����/���1u#�[��3�#*8Bq	���N+ɛ��󺈷[r�x��,%M������Ab<�U
#���tdER�<�i�+L�S����Y�@3�Z�9=kc?2�K@�O*Lba�9	S)��P��VVe6ㆳ�p�C��wd�d7�����Vw͞Ԇ��=1,t�{�����Ԋ"�s��i�A>a*I߉&�A�GJ2�v���&_�@����$��b��A<�"�,@��R��;���l��s�A�&����vK�={��HG#*�>����w��yG�{�R��N͏o�o�vAA�`�wk'H�.��<�T^@�by7��ǅt�d	�e��pf�3:�sl�
��q�3��9�''!�l;�;+V����-!6�z58�;C���DwG�R�����)�ΗW��d��G�;�r�ڃe��+Z�Z�zul��[�Iu�|1i���) �Me��Cg)ȩ�����_�_�ȗ Q�^]Oz[r��2x��C#�1�ț*�Ƚl	��u�{����s�Q�Xa��PmU�$�j�T��(k�����6�ciuc�~j�d�g*�&�J`�B�"���DV�ʄM��+�-v�~����L����;hS�~i�Fs�rF�`X�і*���gj�.�X,��y����1a�鮭�[!8�i4���~�8J��ʨ#��n,�O��o��da@Y�bF�"t.@���y�K_7�ֽb�-�c�s+jX�����,H�*��q��H���O���H����ʳ�	->cM'��O?�=Y$�(L�Ԣ��9�ؙl����b�.��T9ˆ���K��G�O&��$]u����#�'�z�'0�ۚ:���2*�LpV��+�"��=eBbM��k<�|n�ÝZU����a$qf�xZ����E�'p�]�
CS�(��=�X��� aH Q�$�e ���C�w"EcdZ�PF/�P.�{P`^�5�*��%�IS:0PDz]�|�������>�}�[&���n�v�?`���� �G�;7�⁝��K��p '�AO���@�n��
Lҥ��5�!������}K�Y�E�� ��5	�D�%ƣ�*��&&2n^w�j���ߥ��L� jm�"dAt=Qo7�����q+6@w��Y}��B���1e��:Y<P�������HM_Y�.ת���ind�᧏�0H���5��hZ.lf&�"�绸xE�3�T+��dE�����w�70}��/��Mez��3�_��M���8�-�V`\��w|��VH�~��j7S��N�]Y���$)�m�R��RW���F仈h�?
T�8Os�u�y��0��!��*-��$5�6��Ҫ؄9ݿ�;����W���eg �2�9��ѭ<�u'�D��v������[��jmn�_�ز�V������9���ݜ����PΫ�$����-
���՛��_apw�<9c�L���gծ
|�U��u�=��R���6��>�v��z]��R���x~`������'�MI���X��Q�H���GV�Å�/�s4d��l���:�����p��(m��'�kS}ف�Eݍ�&B큒Z#�;��a����N��4߾@$ɹ��?b���Lux�+-3�{9�Țذ/ů�#8İ���f�B#���.�i"�Wr�L
�BG�"{��~�|�蝅_<*ok�[A��Q���\���� �MصQ�����'�����Φ�k=�C�S��Xұ���6Y��*1n3H�~J5q������j�+{)����"�5�j]�q�酺b�
���t���R�kѲy�$��ռr{W���@� �!b%5h��Ӳ��rݜ�L�o�����|��z��K��$F�;W�s���h�O ?j���Ws��D�d�	�a��i���(C͵
�0�0]h�"n��w8ud{]\s�Py��tr���olS���RWV�����J�B���	��_~,6꣱��$�+,!u\V� ���%ⶑ�����f�92[u_�L��E��c-V0>���n��^��w�q���ۅ�j���:���y�đ]�hU�f#i��:�_f��_�$7�8�
y�n~�qy�;i=%��m�gA�N��E����L4��v� ��?�$�	2o�����w�S|�]�WO��þ(�u�)^Cz�����Ao���~���Qx%�ȝ���/�JD���0<�Z1�ƕ��&2Í�������X^�Xw�BO{M�k��gt~Uh�rO�P�)>&�0�|�[����_6��YTv�������/�9��U���%'I���*��0w ��R�����r���)���{�oO��d��|�������P��q���v��H6�#����?9��d�t`wu1��ֹo����0S�G&�G��"��C�T��?��|!�u��8�^#5��J�uu�@��Fk��*�6��s��^��x�ju���R��ڞ~zh��'���!=|Pm����]�#	�W���� Tb�K?PEJ]T` ���己�5�������^ˮ��)m���6�͇���w��w�ӓ5�+wqR�2�m�1���^�����2(��b����}�v�Bq9���5��,�쩐n`���X�[v���'�ٌ��h��Q�'k��٣��@�oN�ź�LSDj��K���o]�\=��h�WУ5#�����au鑹�_>����Oh��ԅ�:0�Z~��z��77�fֲ� �t�6q�BX��XA�P�U�G4Hq��	�há�[/+Zd��C�z2U�(q�]R����
	%N����q��xS�t��<�3�W�;hD���o<z&��2B���>��k�l~>U��e�V���交3��"�/�q�H�W��0�d���y掆�p�\��u m7GM���* g��n�fH����[͆`0�'�n�+��{���h3�7H��"h���5�|	@=�m[��>�'4áS}����5������A4��S��P��m�g�?Ln 2�Ep^�tŅ��pş�⵴rĺ�9��ߟ���w�`m��a'az�p_ّG�ۀ�S�8�e�I2aRB���%�)�����c��C�m�x)"O�8�?��7�'C��؅�C��d�h�Z���4Ln�U'j�[��.P�t��g�JFS��`k�.�'�G_�W
�	�@>�~��`�u+�C�����V�>~�nF2#e�li���xt��^s�/�-4�a>�W^����t�s6Ub%|7X6@:�+�ϩ�i�ܶʳ+���ʖP��9@��w��?Y)d����EEԉ�O�ע����Bys�y�l�S纍"�=�%��v�����_2_�3RHp�4�{D�|
G�^UҔ���S�X���͍��1tUߌ��A�ox[dV��m �Ư����kj�Nnc�`#�=$:��"���ʥ@��A�ӹ�n��M�Q�|�.�ʵ.c����	��<��a�]5�Q7$��.Ȱ�h����g�v-v_C���J�U�4�\L� ���r�8�%Ҏ�y���Ik�ډH��l���M4�}�ۧ9���cu4�����f�a�ʰ P�;��e)��i�^R,Ϲ���cK��f����R&��J����VnF�h��Zl�ZZ��CNC�cʹ"S�?U�P^l!���	������� �2�N��3\��dc����%�s&�{Ёv�E�i����������4�9RaӅj�eO�>�3�l��Cg+
���?qY���z�#���&`:���Q<T	� @Xo���^5f��!�`	4��Ԋ��w`�d�o�L�ݛ%1Ӽͭ�:U���k�d�0�I�
l��.�����7|�v�S (U%;+�Q����	=]��G����[�u`�h���~�����B۷�>K��h�[��%2 u����/[hA������B���N'b�����*��J+��v?;�tNРm>W����V�-U���h����P,B�3|-��k�@�=�ER-��Q�j�K���2�$X�
��+�ٸ}c���f��T��O�:�����6J���KZ�`[OXA��}��>K�S>`Ȼ�:��)1�F�_��w��o�emk�T���k2�U��,�P
��q�a��O���qb,g��ע2�{�b��2��C���]����"�s
���S-(�=�(;|D�?�2e\0�X<2�A4T��>���E�b��M�
Ԍx�g��~�ũJ��vP90�9��h�j�6S�]���@4�j#��g���DCdlC�j}���T�I�Q��������1=϶Z?C�զ4��4�3 �2�PcF���c���Sr���닢�ی��*���q�s��gxG��4eʯ�9���=M%��L��)"=2�-�z�HX˦& V�������A.�s�Jn(�6�=��p��[�/6J�.]��G�)Q'�"�8z����ս��w�cL�M*�Q˞,L�2�P�R�H�\B��"2�n�� 7��2��I&6B0����7�y�
�B���_���1ծ�⻜'\p�.�C���"����ˍL��i���s?�lVy��陆�ʞɓ�jS����.Ч3�Kqd�<:OzQm�f���%��v��4��w���"v|�����˾QGk,T��ˋ�7K�����=�z�l�c��l	�^��ɕ���+��$V�wr�C�8�"9�(�}}fu+?��*`�Ux|��a).D�o
r�E����ع)�������7p��a/e�Ɨ2��O��%��k�!����1W��
p����I�9䄟P�~���TO �{��K=�����m��Q�,0ܼ:�����B���=����;v����m7��]0�lA j�&�3�=n�.0����$��,��:�j���k���,sb12~�Z�ϲ�`�(�>C8�W��C�����V�LX�
�Fw�'\1�a14"osfA1i�gU��h�dE�Ȝ�W"'v՟&ܱ���Ӆ%�^n,��ơ�?�o�6.;�鷞���uP2�=���2j��a6��Ii�$ͣѶ²�$T�r�@��u��J���"��M�¦��?���I��1��\޽����d&�k?%Q1��n�(�9�Y�����bp;�U��_��*��v-DED���ωc�nB��:\�C=��?�⃇nssX���������vr��Q�t�y��+�o�f�p�Q�	9#�"z��U8��՘b�{��
�Ga�]���]q�����eq��0\���эXd�=�?D�J�vc]W!&����V�Ǵ��p�{p5x�I@
� I,L˯�������z�|?��n�gX����,|��5��Jq9Yʷg�)��	���fg ��z=�$P0�j����;��2��c�)T��3[6~hZ	�(-XKs�e~���}*l�����Y�I襔�p�K�Z ��X��:^ n�P����l6-'����
�.�<���}�����t�[BF2�x�x`}��C��bu��A��
e���$c�$NΔ4#x�T��
���F���y|>]���`0vxZ$�o����pP ��>�흄Ȟ�4mK~ڶ�Fj��U?d�����"2��1rD�z��3��:	�����zr/\(�J8g�a��2w��n��?�h|�)�����݆�Q�E�M���D4����VkX���pnf�Őh����,R"R; F����.ljX�i�����Np敲��|�".���9*�/uD��fp49?�,K�s*5��x��:3R���e61���r'HЋ�_L���M�z�)3����Ҹ�_�S\����I@���X��YoOv8��粶%����,X��?���x���;�Gk3�I4>�_9���H�7AmdB̅ol��6��X��lY.���ٔ?�|TBP+�q�uͩ��J(�Ij�t��GW���B����3��~��A�{.���ŋ ڳ���=˻J�YA�C�&�u6f��!kn�O���_,-͠��C~I>�7k2��Q�	�d��h�U��/�܈�R��>�%,�*���4�D;J�|f����k���@��A�|H�"�x�h�5��MƔL�j�xO&�!}��%�(%?*kX�5�b��Z�v�OgΈW@�V�{2�t�Y��b!|����N*��%<��[>,;� ��#E��iX�=S~���=7�^��n�OS�Q�Q�+��3I�;�b���gLH�vRJ��{t+��NO�]��d2���`�ᠴ����+��Q	pFbO�D��PM���0�(�D;��2]m�:�Q!�!���Z\�;����=<�˖;��\�c�򧀈Iv��`�K���2X�ɴ�����z
��aG�t��ᴂ�۪re�u�
�Q��䒲x&t]b��Շm)�_��nn��m���B���8�`1�B�a�kIѝz�l�͘��ʐ�R�m�]u�Lq!����~ɝp�#e�A�5%}��.U5���)�	s�1I���s e�Ⱥaª_�jΟQ
�ͪ��YW��I6��֩ƭ�@��W�,����� ��<ub,&iP:6*�.�1��R�c�=;�sc�(�G�n��U-7�Y��p��� �tא����<��dl�ն&z����[�b����9���P զ']��)��C��c�� w?�L��\��9���y��ɾvV1I��,�����(ր����?�분�T�T)]쀝�?��3���P+t�f�� ��J��a�P�0���aP�m֐7�"���SV0��ʊ�;�k�L�w���c@A���<SY�,�z��_���P�~�2���iB�*�h�w*<���2�J�T�%� z�~��Lؖ��և@�yt"�a�X��G5��A��ѣ�F���.��o:��J��r���xxͬ9�i>OKC���#�-�%y��O�T�LPZ��%j���|���;�_E��A�8�+M9�m<���j�٣ pL8�w�C|����j������"��[y���eQ70	���4:���n�$ľ��i'0���9��,-jL3^����` 4 ��)�����fhCo{z��K��(�>��{��0F�3�έ�%���:�Y�:�"!�7��`O�0��&>��� �c�8�������&�DN�ĈڃITA��I�����B�=H��ȫ������k�<^^�#b��_���m!��'�|G�N���Nx��57&T%�X�V�����ic�F�����"҈�u��;Rb�X�V~��х�g���ى��?c˪q�U�l����>�'Zh�=�R��߶z��Tٺ��$w�oE#v��ҫ8Ql�4r��Y�>E��T���B݂��#@�j�rJ"�`���]W��~�\7���2���H��1��t+����Ր:��n��㗮��L��T�;�p$�5���~�S�)_��S��3��@q�8��j�QkD��P&I϶����9�'�O�E��M�#E,`�gڧC�a�+�*&ࢋ�2=���n���A����p���.��{��1Giq�Rق6��e~}k�t�]��1(���F;1E�13Y�'���i���.q�����9ť?sT�B_�l�Lp�ڢ��D/x���F�]
�N�\1y�q�����
y)�;�5�e�x4�L�C����C09 /�6}M
�� �1%�������[�SEBX�e�DrL~/��/C��)����&.nIH�0bt	K�:��3��A�&-����y�|�Y�)���1ļT��z��B�n�29��_�z�v[���إ�*-n'(��׮<���y�<<σ�78_k5w����x��Q���n���Tdm�\�6`�БWH�V�=$�fdGQOÃ�C 8�Jή��p�s	���?&�Т���$yD�'�iM�p߳�h�`�g����ӣ~Wc��wB������sM���4MЇ��g�x��Ag�z�i@ˤ����H��A����n����V[]����j=8�s���V3�T1�]K��B��1�v�������+Vy�o��Z�>\���:��۝I�D�*�B�N� �>��od�U�1	�����2��v�kZ_O3�A�Eݣ�wlk��,����Z�����ڛ�t���ˈ�2�?n��g#�%v�(����Ŗ�V3�'h��W_ �8�ڃ�v-O9�w�իTA��������Hl�ز�y�����x��jQ�:&�  3	C�.شoT��i|m�i�|��P0��Z�K��Ұ8�F`��a�j���Q?e^�Յ+F$=C��2^=�c`	��>�X嬚��͠[��q�wb����2�|0�P9y�7C{��C"�����7�!%c������D�K����q��a��Pm������u��cP�x@Tn�)pR���^�i~�^F7�T���cTA��f����a��q�,���K֔��8�V�ʨ��xxԚ����4�}�f�
DvUȷtHz��9b5�h��H{7H�V�>�M@�@��S]��Gs�{��"7���B�a�aj�xp4ݐ�+��r3����˱(�I������:�fa��#̧�2��o
��I���ʝ����j�6'W@��=�l�� :1m���	�E�~�[.�{��l��r�B�>#�����`�t��L���u��_} ��	jq�������=_R.��{X���m&`9��w!Hl�Dk��l�fa.10�^��=j��sp��a���`��\��Pk�:��'�B�|&�'�d*	���΀������m�����zZ��_�n�^�Y�+���ȵZ�ܳ'b���u�;XRR�O�\�h�`f�	�V3^�0��z�t�i�#�;�>P4N{�w��]ڊ���/�B��V�~�-�nR$���e��+M�4��8���k�,[�MВ�a�``�m]�����8��g�l�F���ǟ�Y5 �UlmB�ܠ&{�Ne��X�4�C!�M������EKb�.tTMRx��õG��<�ܟ��v�~��g�z�x-�/ɗ�=2�6��Eqx�z���ze�{ }�����ɺ���~(�i���/9����|�Y� �Ņ+��Z{��0�X���X����,b��(4Q�Ϊ������a.T��넝��R���#�pr*(8�((
��Y߯�_dD�d�߿�+{)����OI��`��ma�o� JK�b�68��SV���O����+ �^�uD��U�ٸDr�� o�%YWv��o�����8��^���3x�qbsK C�b[��TЅF���ݒ6[P� r�kš-�X�ᅒ���������3�K�wRq��yS瓵��U���dI�V]�R|�j@�x�s�� �k}���ǤВ�e/��K8���܏���ڬ`�"D(Զ��S
��|�j�q�g�f�2ly�@���\�)��=[�T��f6���7R�p�����X}A��-_?�.�¥j$
��@����;C�p�W��,>���<!�2����>�$Q��5�#�>�����?���%#]�o���:�:�GhY�~J� ��o[Onw����'o>/��F�Zx�^�E��̽�o2��D�}>�Wx�Z5�ޮ�W��`�U���KUtl�mn�L��ݬ�-�;0�ؐ�����cJ����:Ʋ��G��+�0��@d���֜gV}5���� �����,8�bczs��ׯ�o��ŝg� E�Ȥ�
�,<,��kK<��Ut���T ��#�B< �g]�� ���S;����ލ��Q��Ǧ��|Z��[�3c�O�5�l�tH_�C��УVM4`W�+_��O3��$X�M�m���tqH���g���gXc���qX�,_4��p��]6
����!{�ȟ�xm�0�Z5h^��g��>VF.�٠�{z��P`Mc6n�^=��q]�i$O?,Y�+?�vh��a�$؈�}A�,W�O�ޤ�^�S��{��11R\�:��XZ�
�����[�>�mr:2oТ^��	�D��W ._�-^����$�����區C����E��+��,�=ϡt���~��ϻ=��V�)j��}�,@�	�HN~.�c^�x�`pS����]��Oc�]ʤ�?�	Wl������N|�-�L�3w��)k���H� Q�a��c?1��������	ی�ZN�ʿ&��"��཈*u���ia�AP���O�ѱ0�ϔ%��2��	qm$3w���6o��R�R�3V������� %s��Hwij�X�;/�K�IF��>�d�e�a�;Օ���U����3���H�Π"��1�()���A�L�����?M��U5v��V.�k	��7֬����J	2.�v�7�.㼈��v8����7pi�T}D\��]�4�������[ɿFK�o�Q�~��1QV(���@/�;�{{�#�b ^��r�qW�٢��+������X�6����4���j��#��
f�b�Y���D�MēS8pA�)�
Z2EI�fV�������"g�H2�v% 6%Þ'v>��*�l9��+?��\�3;RI���:���/ �/G��u�F=����|�PS \��)������{F�i�ٖ߬�G��mcCiD�P��=�p�LcO*��w֩����ޅ��a�Z"(a�RM7�H���J	�p��l����+R;����ە��Ɇq��O�Z�G��� =��E}��Mښ�(�o.�ܰ�A�1nST�d~S�+o�
�Ħ��uYp�.M�"�8�]	.��ďzr�8s�v)�ne��F���
��,�Yꆴ�R^g -)��{B�g�=�]"���g��������Tm	�(	kO�҂�Э���g�&�|�>�iJ��t��"���x JKЪ�k�RZ��/ݷ���!�����W����8���������F��=k�=���MJ����NIx������J���ďY�=t���������s�։��|6���
��L_:,XM�[6���`4A������	�~�"U�䣻7�E
���l�{�h�e�sZeĲ�|���W�E���`62��㑝$�H@V$Y�/_�а}j�!�K�0	<�Nұ'm��7�p�������:���eM��Q�c5�ǰ�&��L�w���؛�5x�(��9�ǭ��V�+(�dZ"�b�t^yK$,#�M3�L�X�f\�L;����WKB�:!BCBa{��P�\�g�N�i�;+��ߤ�:�?�56zً���4��[�A�~�p�z2���g,�g��o]m��6����.M�y���Pn<,$z�����s�$j�B1l�&���?��7���S�rJ7aql�
�7c�y-;�$~�ͻ�Չ@I?�� ���ĤH���y����.�4°�Ǒ�!i)�Ǒ�.���b�jv.�m��5��<���,�H�iL�{����p�����.��I�Wu.�V�AmH��R�қ����?�=E'���
���&B�h�a���+
-�nC-l��o��Uϫ���Kx,�1�q�F�ҏj�=���U��Ч9�DɯU�d4"}r�>�/ȐvR0,m�+�EEz]ڣ������������kйПy��L������k��V�ttLl��zV��߆��m��S?�t��ЈUz��7Q�p�8���^��4�0Ʉ�p	]h��LIb�$�+�������Vk������6��R�m{�\y�./g���g��s���Lэ}�Uoe)P+hA��~�:9أ\�l����7�)�P>�����p۫?�%z×� �p�k��|yg8Z}�n ?|�g ��3����O������&
��}f�-Xs�Q��-�&it�p�~�Ix
Ya�q��i���ڇ�HpX�$��~��v�|K�$W.��s�|?�θ���ݫ0ݘ��E�<X�t���3<1���s��lQ7LU(;x��O<��e$�S�m�o�6b����L��3�ȯ�5���ռw�x¯5JdL6v�����:C�t��ݒ1�֡8�f�*1в���[�Q#�������,�T�((��o��H\��ɋfK��V���rx�)��̏f�Wu�9'�y�.�5J�'���P�z����"H85o��Kt"YО�<�zO�J���雞��I�٭�W������9^����1�**U$��8u7b<ۀr{s�n{qT�ߐ�b��b���l"�@�R�Z磕0��X�r�D���\��v��}S�`�!7ŷ���θ�KȖM��#�ZeH�R���>6IW���r�ㅮ+�ԓ�ۗ���'uy��� ��y�D_@8p��7������[
����I.�C��B�A��� ��,Jui�h�B9�p��Q��M�Fa)�V��Z�0�P�j�:zȐ�]Kܑ.Q֫���V��J F�Ē�&�Ӱ�#}��s�q�^ ���-\n�q7��%U5|�=�w`��rt��@:&���S��2j�7B�� �W�:��M���Z�r��j�1��X�jS��Si!�o*�&�6�W ��[�RKecJ��;�9*"D ��	?�У��)�V�j����*�w��]�/�J�y�M˹ԋ���3D:īQz]�|��S�e�vK4)p�Wdi������U�$!�wLQ]{	�5��c���_���k���̇M���O:_gg��Џ}5r� |�@�XӛΣr�p̾zݾ�#�F�=������߿6,ΪN\5Sm�?�q!1-"�};���I��P[�"~sTȝj�3��@�������QKwc��5��0�z=`K!:*C>=t�j^j�hJ�����ɽ٩o>I��X`>(�4�b����h�{�vz9������P'�=l}ݛ�sN�r�Wj��.�b�ےI��C�Y�`� u4E��w�1A�1fb��+�8��QƮ9��u�6�D�(��KjH-����HDr6K��`�߮�Yٟ�,5Et֫�v��'Y����^�1 w���X��t
4N}"��d��m4�Ky�9�L�+$�;5;��/�?8:G�2��5@�������wT��H���kU��!���̀����*�6�@��2�"~�a�nOr��w:�أ翭��t�1��,�g5p��T�(����/���""��}��[�XP��%v@,7&�D?�?�=t%$zтk�fZ����΢�e�ʬ/F:r�����4=k��(�S�p΀v���84�w9c�4��Y��1�$�ۂ
�q�(�NMT�|���B-�R�F��S��O��r�=x���-Ļ��v,6:��#lv�1�A[���.�݆Wгf�3H[� x7,�� ^�*��q�3nf�Ă8�yQ>D�.��� ��RI8ؒ�I��T�4~��P������(5x�ȧ�� m1��+y�'��f��������ɂ�+����0�IEN�x����~A��?`˴���޹��TE��%�Uz��[�Q]�����Q/p@�G��FU��������.��z_Q/�~��Pٮ���r�����[���B�0y��W�¸�{$X|�=�@�$�P�5�uE��ʹ5g��"7��:a����
�L�A1"��Y�hb�9���sW��A&a[�����ֹ3=�"c	�S�[C���s�\��vSꗟ7�ďp�`�z��`1�L>5_����m�(���lĽ��:�Y#�\�&^�վ��ևӢ|���p���.�mM�qg�Vi"�h����罗,9ٸ�(���4m��j���v�I���,@_�����g�%ۚ�"�Z�3xq���cC���݉�������4U�ܢ-Z�Чέ��+���nV弜���f��bQoz(Wm�y�s�Oy�)kV<�Z7w�,��W�g !�K��;��� a��g��	o@�V,�V�_)������7V��.�z]Z\�V��#L�ֆx��]�6�Q��� *�r�d��؎�����a��Y�?m�� � �>7�à�g�L�?�B܍u~������h�v!�
���53��0v)�نf�N2��j?@z7��L9�fY{6 �'�����iq7�Z�������D�>�Nf�-���PqL�B1	��O���-�I�x��vW{y����^�[('�Dd�^���L����LV1�
�Xr(0@2�DyԹ�3�n��;/3���`h���� ����X{e�M���j0�䊰?�fg�u)��cC���~UFyI��R����I�ٱKY��"Y~@o����&��+'XVb���B�qT�$A{+�;D\�:ϡ	V�R:�O���Uh`<�v99�z3k�5Z~�Tb�z���%�;^MgN\��R+�w����]f!�9���?P
=� �-��w�W|��Q��:y�Tc3p����d��q�>`�v�k�	�3֜U���k���:�<0-íϿ�HVo`rD�F�KPG�-T;�.�}���T�60�s�?Ynl�=8�j<̀��9b4۟/yڞ�A/���X�q�ն�n3Bk= $��g�u`3x*O4�d�Q�`���2@��&��D0`2U���}I�Nv$\y;�F�J����	�S�>z�)�ɔ�ǌ�X�e��V�	1���T0و=�����	�*V�]��9u��s���]|�<���ـ���7@��y��ǟ���~��������.^s���0��aҙrkhX���wL`i�����/����!}/������z/.\�.�B[�8�/�pT�E9��Jއ��Þ��dc���h�c����
����}�p�� ����J�aȂ"B`��7��1�R�b?`��~n��3�@�����r�����9L�yV�d�~�A2Q)���YOyZ�"�޶�Nб8���ՊYf����Vz���!��g@���P?Y#MN����Afu�C�1�!q�$�yࢠDTo���_x0C�݆��!�1����k���@	E�#W%����{􆪆~�njt��U q�}������p��*3�t�M"h�}���_>>�C�\��JZ�8H���� :P�Xc�:X����s�V��q1�X5�EW��F�R-%{m���:\kV�K�7�И2�nhߙ��a4T�=Ϥ v�3��7�⇫u��؀�~���'�����n���x�M�J��F#x�4!楖��@:b'����8&���V(3����'3=��K�b��}7������l����Ǉ }\�L������B��4�!�����?��d��Jj�fT~e?�%���j1ȧ)��8:#Q>��p+��y� )
39�7��w*�7N�^�2�7��xNe�iu_�E��۷
u�O]2��˨�,�^����-�>����3#;�~����iE�zI��$e���2��C�
�G7�6�K�h���B�����0>/�kz18�<JR3�����G���,L}�1�ߞ���[����w�NV$mJϿ��n��U���}@v=����G��cq�p�USX�z{f��3��QC��q{{�P��K���ƍW��z�e�v#�Pw$+m {�4�(}���BD�����x#��N^2�+�ߴ�wD�7BwX>�R�ym�j�!GR)����B\U9�m�	�?��������3*��C<e�p�Q:`v��"}6�x��t�����X����)����U�z�<��B���?/��Y���[f�̟������x�u��I\<�$v��B�	.�=<�����}��7i�i���XTq�p���Arωq���P9���΢x=W=c��t�yS;��j���Eni� �MvB�'Z�!�F��������_�@@ڶtW��K����Գ�h"a�B��S{�E	�~��[4��:��ieq��<�|H�"I�@��^��p�c�Kt�{y��[LW/����y8� S���y�vl�u����;�:��O��P�����~��ϐ�?-HQc �u.��s婢�(|���i� o�Fp9.�⿫y�v��d�<7���Y���^[��gl�W$���J��Q�Q���<�-&Z�VO���x��ݨڢ���Z�Q@d��W�����-��oi�y4�a�c�KW�Ÿ6��5���,��K������+�rS�=�)�:�s��x�lm����g�|w�,I�=���7���w��Y3di4�r5�rF�.O[�FP*���pLV(�����9�p� a�� �NV.�ai�jL9�o�����͒��'kQ������'ka(Ӻ�Pj��B���8�s��C`��� L{��ǗJv+膗>b��VVKO�%���v���|���G��R��n��H���8a�/�X���@"��=9xo��X�����*O��n�7~,�n:�V���_3NOFmڙ��h&#]Ѭ�C�_$&��3��t��},��G2���W�~�Y���;��[�T;�Fʻf`��f?�]}�3-�x7�*����jR�W�~�����4��l�()PN.R�9[�+�`ϱ}*���]����^���jb?w��@].��Kw�گ��A��F-:X*B�pz�D�0��E�;��d�A�h3�X��dR<^v$��3ʑ܃�������E�c��4,v�97���WH���4��Vs���p7]T��bM��+R������[_gčM@�]�{7+��4�»k��r5��L2Ԗ�&3d?�@y�F��H�6]�����u��#�
8S�����&� :_%���-��H��Y_�V�(Y��/`�!�:EFa�!�`&���, f������P��|�i��4I��*����,�7��WB�	��y�ȓS]i]�;��1�xԷ�T�huxf]�ژjmQ�I{w�PB��e
�ta�YQ���E����	�yr���	�c�r�Z���R��ב|\+�����!��F ʟ��B��r�q�%�_�	�px*��8���V@ES�-׻��*�7������L:�X����	\�}3Ng9Zgi8l��R�g�U��-5�Φ���Q�(Wq�
�Ѯ�+�8��g�:xB��VbE��\_��8[�&�C|U4����L����Τ��q:WX`���蓔U�tS3��B-��G&��]�Dq&�1�5Y�քo�!	�����<����,�>ywDh�3��k�d0��C7f:��>ltν7�1�Q�8T<7K܋ʹ	�P�K{�лBm�m������Q�yxl�9���G�!�jEJ/�f�3g b�iҗ��7��s>;��_�Y1�Y�����6z���(a��Й]Ę�wM.�L N����*����Cha���2�K�֬� �3]X�&�����(,��	�4��J|�<\�6�[�r�V��a��b���=���4���b�1ץ(�ji?�ݼ|�4�;�Q��tQ��!��t�/iz��9�`-��B~C�{����[B�����˩���j_ ��~q��ؠ�۬U~��iGVw.&mF6_�,�`�6��T؞�t�e��ߦ�cбb�4�?D�� �����8=�����^��&!�F�Ji���.�>�m3x���F�&d9@$/d'�fټCG�+nB7w�",9�g���$�h q#'��!�RVc�:Q�1ґ�HDaW�x̶�D&&R@��z[�T!D���8���a�G���ۧ��)Ir出I�k��2'R�����Ns��t !�02d���ADBhr˻�g Ya5��}�e��U
W䷋X�I� �3.6�c�6vk������O�Q"2t�(���(�B��	E;
x�YY�Y����i��פ,�� h�I(25���]�ѫ-�T@��LcS�W�����Z����T�$�K�n��I j�{O��ǀ]ҷu�ֽ�)�/9��}��e����9k��X3Z����냹]D���m���?s�uP� s�P㩜�W(�֤Wc�Y�I
����":���R8��Ј#�ʘqY�Ӗ�&��h�5++ӭ�ϸ�J�JT)!$�C��տh��L�=���&��V������jBR/BÓAb(�$�؃>�j��z�Y�u9N!�D��&��������M�>�+x�Z8T���T�
�bk �䏊��F�[��Wj�H�pq�}�PCȏz���$��3�#j��݁t�]�4�6T����N��Aj[��װ0��B�Ƅ�l�4�Z�fO�[A�,z���#[A� yltG��nW�NP�>+���]�����F�+�q�|H�����R����AfN�1,R�' k��9�~��ޣ��0���
�]��
�5j2����䒠��֞6����T����m>�&��q�i��S�����ꤍ�Q<�)�Ŕ��>I���շ}*R#��m]G#�z�d��$��d��];�	$Q�>=���r��Ŷx7;�ۆ
���Ed��8I����g�\�i�u�F/ _�������/�אd]g�.(ZB��9��ҷ(U<�Vr1���z�/ߞJ\�y8�:��u���o�Ԉ6�dF}�m��it���z#E ɢU������MAl�(U4�=�ەBh1"q�lvd{�s�1��R�/�л1u��S�����S�Y�r���C,�L���7Ӎ��ʷ�e�=������;M ��^�(]֊D0������@�\���B�_��}!��/����K�ASݯ�ǷjY�;�H�:uR[gyɗR6��#���z�<�qH��$**��:���m���$s4�j"a����jg9��,�;�~G_�qD�a������ѨBqQ�l��X^&����}�]�6H6��X�n�=}�B���X�8
~u�q���3Co���,}�6���_6��w�~J'^��ILku�N8+?P�v�Ҡ\�_�,ٽ(G�ܷ��  ug��.Iu|k~�C�ӯ�f�ڷ�l���>�a��//\4�/�<�AA̡�݄I�4��c~���я�8z$�-%����gs����E��,<m^��nPP0ck���ߊb:D aސۓ�ĎI�v[�XGr�b�Nw.M.���c(�c�����9���b6�4�{E��s��h��d*R��L��\C�������n���ǌ����2ԇ�9-��Ib����J��1�ҊԾc�M�"���ч��iBR�x�Cx���,���2�U #�>F(�g�(kW���K<�� ر���8�����E��1;�&�y�������6�N����"�I8�2��>S���ůa��8c����|o�dBN��|�ΏH����?��L��ty]>_v�5
�g�G�a6kjp��9��1���aGyr�A<��e��p�o[��#�Ƃ���'f�9� ��1z^]�.�p�F1�MPDS�ubHƒ��5��D��(n+u�l\4sO�c���\@F(�ř(y��,q�J�?��j]�X� {g���qE���s�����h,�8���^g$��VH|#�]PQ�O;�5��'5�tg�S�F�Z|�U~M5�H,�oM5)�@���x����a��aFH8V'�u*�5%�r�^��X3)�'o�}��*x�5G��vIgF�7
���e��|��|�]��D���{���������S���
�D�n
+
��{��@?M;��up�xަD?��x�~�el!�wc��Q�p%�����������6�ʧ�	�)�����������K�R�ڕ��`1W�8�����XUEd��T}�(�eV���	(6��k5���j������_c?u���Ҥ��a_OBu�,_�ћ,�d�����QHe�%B�����G7J��>tE1Þ��/����WN�
�Ix��9�3�1^�;Ə�u��]�_��me>��n]�;y��x�ކ��ȣ��M�m��>���TQ��װ.�y��|���j�e0+7���)��T:.�؎G=%��s�X�BF=˞]�n�)7	1vy��J�����әJy��f�J��\�2d?^%�@џ��)%s�65<��v���?.�}��[���,�[NP�8�)���R�|��T,��E��g�Q	�'n����ltEү�
˞?�h��,���t��j����2��6��Y9ᆐB�ܐ�n���N���,�!= ����w�0k.�B��:��ŷ׍���	���E��I�����r ڎ;BM�bc��6���IQ9=_vjC��[�g$e����t#6�i>�vL��s��Fy�Z��I��tLM�4��g��M"U�?T����[�n}+�>������׼ZK��*�A��f
A)W�jFA)-�T�w�Yx;�q�kN�{eY��\�|���%T����������~V�Q�W؅�G����_�Pe��ZV�������|��~M�e�iF��]r�v�O��A�U�i�Lk�[�Djp�]@�EїJt �5d���)���YOK�:Mt�I�g�o�RD�fd�) �i/��|��-e�*G�˃H�:DYc�A2�����|��	@�3�;JC������7��$��QR�vbJ�n\����л2��m�q�J�-����#��'2��cJH�b��WJJ��ӋU�|�\GN!��Tʲ	 \��HS{��ȂM����8Tz/��Np=k�V2��{[
��C8Y�e������WR���J~����� ���@�E*:�R�M3��V0#�� ���������(a�5ŗ��倏��u�@�|ACYט/����N��\���=��/���l<���<%}��3�O��/eh�cZG��Ħ؏�d��-��\��J}�\�:-0P�֠sw��Σ�r2�㆘0XH�{B�~^��a���4�Qf�N2���t�$��&ϟ`��"lȶ����*����I��kt����5&k��c�﫱���6�Z��5c�}IT%��-�h�ˁ�����ވ�����*�K$.
)�t�B���������/Ab���)N:�8�<T�_���x�dTh�)�pΙ�'b9O�}�H��X��h6���X�ݐ��6iE�� �N�Cn���"������S�;c;���A�>#�F49�}�αR�=b�ʃ����h��!�q�ҍ�(�1����&c�&i�1em�W�m�}��8V!NN���ź�!%a�)��G�8�|��������"���nq�Q�y(�	4�p��w{O�QG	�j��lk�4����������w�5k��9�{,���~�9����W������эԄ��?�v��kr򽫾=L֋
%*u�P�[��R�,f9q����f�^���P���1�����K�S"����S�u��G���Vjp�7���㾗3�n������է3q�n=Z�D��7D^�U�0Í2��A�W�!��3��j��������e0�b~b�*B�H��QH�B�!�Ӛwa׭,����~q6u������� yT�
��7�ѣ���oe�N���ꞏ�
8q�c"J5�aHuO4�?E:��R7��Q���2��=Ȋ�<[`,Z�T�8�o����mF�:��	~Cy�H��8�F���?�_Jm��b���E���^���S��HߺD'SΞ��"ʇe�ׇA|:�e9��1Q�ɡ� ��4<�g�#�W��+�lp����D�e�4n����bʃ=��b%=`�vX�1���'�T��u�#�Q�$du��E� ��X�f�I��Ӗ����9;���o�.���'\�6s�wr���v��_Dd:+? �mD�6�S����~HQz�eP�hb�C�B��:�y[�1T����n	v�!^�.��ƀ��J<b�T2����OӸ�]K5>�:#9�t�q�mX��p�A����Й���Vn�-��[+��v>��2��p{T."� w��Q6�"���A�X����wO�{DƈE&���㥓zI���;$2����3��'m�5��UҘ۾D�mXT�e�����}
�܈u�J�����"�/ݼ����P��	�H�lz�&�1 $=p�A �#0)�K5[s�P/�e�U0��<l���ޫ��d�k��9��V�~h����gc4����ٹ�& -��}tk|�����\�$}'�w@y��L%"k;�g�V�^.��PY*8{�l��[M	&�P3�|>����%�N�o>J�By� �7� ��Ѩ�S��Sbέ؏����`�z![vz�+�������\~M/�7��Ѐq�����
�֙��r�'�z�F'��l�����v4~���$}����/�j�d�~�o�6B[�]�� \�`��H?�=I.k=��DuP��;�s��Ԓ5��ƚ0�#]��g(Գ`�b���ѺU:�Vb#'�e�J����t��|'@�g�������hR�@����k�N�0Ŕ���żH�ʝ�h�A�s�.4���M��basp����f�����\�F����@����BT�Ȟ�&��E���4�\L�\�i�q�f2D7򤕳����׹����qy.TG�D� 4.*�N�2>e��	����f=^V)�K������=Sm1
̲��%���]�^���0�=[\�e����^��6O=�3L�r'ΑbwӍ�>��T Z���
ղ�Ѧ-�z�/������s�2�yQ���'S� ��&D�9+ �4z��k�N��](��|��@�Nm2
��j�o&�-�⽟g0e��S�Z���8�n�E`�.G9C=޶s��!��n�>5e�4�*_��U�61����Q@X�te �HLCccӧ�d"̌�"7�^��[@�\	0�ܷ�8��N��0	�Nvv;�"���L�)
w��n�����Oflp�t�TvJ
;e�`X�Ժ zlt��i)�������ު���ʷIV.�zU��������=q���)�����x6��#�鴻�����@3�&��YV��j�8\�&xd(��V��5�ƛr��ꗱ�3�_r�yi�VI\��f{
�Ar丢G��3���yP���WS�^�؇�U����1m�i^���G@7��k���5����Ĵ��9��X�p��!kF0 �e{�M].�Ӵ���s�'�f������d��!�?�z��Px�7u�p�`��_hH��O�hͧ<���Ȉ�
v&�����W���S�,��~�lI7#2im�Ӝ	��F(���p
�ψe/R��G$��<2��+��1"�Z"���{�3��%@�v`�
ݲu�x�/>\rҐ������?�"���a1���;ٯȋ��+�OymL��C�Hbr�����"����刲����Xq	 �s:i�.$�姤
8��륮Na�YYFQrw�TB�T/�����.�'YN{����O�}kdS�ZR i�Z���a�*��42�v�G���%�Ji[|Df�()s�s�m�"� Q>�%�g�����+�Oi/�8���YWav~�+������.�'���K���v�>���:�/̢A\�j9�,�	����q͗�#7����\*O��&x�$��4��L�pe�PL�k��0&����d�К�[r��	j�R��щ�����}��Xzb��C������I��"���.Y`gw
ZyI�`8��[�x��� ����U-�?{���?�M�lLsF�y"�*�&,���A](����6�>��/v�RO�K�N���ݏwR�#��<�D�����!?��P�6.��sv&��c��;	����_ ɪw��g
_6[��I����^ߐ6K�a7B$���,4솼|
|�˕ ����X+��Mv�r&��3e���x@t�V%c�K����m��a��n;(��>�\a��cL��Y1�N1�I>jkf�	�KG �\;�q�B"�Aw�4��PƳd�nG*]��A{7�پ��\4�k�}��q��uW^��� ��w���sŃ��B(-�?�Ş��-��@3�Nti<�}���G�<6`��UΞ:,�1��V/:��P�Y�S��,W��������?���)�p9���Č��q<5	ΦZ �k��rZ-^^��6��2xTx�/� ��hgjMf��Yj	�t ��9�����"o-�"�L-�7`b�W� I�Si�&`A��"��,]p��&�Qkl|����a�L�ž��(�B�,FF:�܌��%�J�f��z;Ȯ�m3��N��ܛ�;��hQE��#�(�"����L	�f���;�g)�$�2vH��Jh��͙UBņY�l�وHF����X��[+��<���U��"f�tC�����cj��)�;�.�x��I�Z�̳�=�޵��N܇��ԩ1j]�Px�Yɓ8���^_:u�v��@�Hx�Y�GƼ3���1� B�� �ʔ�������x,��r�EV�2D����{Y�,3��݂��~��l���$@3X��Y�
<�1�2��]��b�!"���v��m�/U�Z�3#�u�}�@���*N��W�A�����&5�p�/^�����G�6;a�9���CX�wL;C7�#(ЁZ�8:��A;% �u����h�S,����Y���~<����"�����Ҏ�W�}<��}e0��o�:���C�)z����2���?�������5a��4�3��O���S�5�n����i^ڈ{D�	4H��!�Q5�&��~O��6L��n�rJ߶QZƌ�t}t�?�rjf��ͅ�/~��2���ĨXl�~M"���Yo`}:{��S�oCh�'Dp��@Уn>��n������A����X8��Nu/�1�j^�5�x�\]x27�l:�b�X���_�66���%�A���'���(��R��0���*�A�_�fk�2lQu֜L�ʾ�+��;'�>��y�߫ ʰ��`�c����ܩ����}�i_7_ߴ��vĩ$_/�*����T���= ����?���^:"���ٖވAܡ�!�zA���W�ey��f`�S蔑�߿r��=�h�9u �H9=Y�)o=c;\�b*`�����6��s���3�`L��D�# �?x�D�4R�Kv�c�Q�1n;aK�F�~$;�TT��F�+9��0%p~Yf�5L��ٶ*�ަ� D/�e����8ް���f����{��µ ����S�����a��'�G4��NtQ�5�h��GI��0�4)�Aq���uN��B����Eb�P�}T��ײ���E�W5�|��+P�y��U�.�?��?��=����0�U�Qo������?|rǣ�Y�dE�_����-���K� ��¨6�#�G$����i�p�'֊?���6�\F�N"6�yD�JօOJTT��H3"_zZ�Y�<�mI�i0|�V��q��(����v��?���f0mL�V&tu�<	n=�>i���� G�zYD�r�*�i<�I����:��	6�q�G�4��/p���zQ�,~f���UvH�
���:�̮��I�	�Vm��e�������f�\�BF�7�� �� ��O�#Ƃ���5p�ߩ��<5h���PE�oP}�)��J�삉���l>\��Z�mJ���
M$r�j�"�-b�9�A�j����O� �ھa��_�|iA7�'�:�0!��0f��Û'CɄO)��=�+v���	Ӌ���K�>+F2�yE�o���U*]�ɖ��Jx�i*����P�0Q&/�pV������|��.N�槿�{���}��C.��ߔ���M=D4��F��hm�+�՗h���A��G8��}@H��S^����s�[c:K_}d�����|Z
/ƞQ􀚺�F}�R�b��pwa��j�R*ݲY�Gcj����P��Fk=�7��Fپ�vy/?_�u���A]�n� ��u�!qt?����\L_j&�:V%�Z�M��Ғ44<��tb�I�k�7�1.��]2�.�Q��*dH�`P%?�_�ȣ �������m�`/e��Ջ�2��n��S[<�G׾Q�b��E�m��SF�{�Ʈ=���`��W��ө}M"�$\)}�'���e�};�މ��:��C^&���q�A,9Z"�Pz���2����b�A���pBb
s9�^��Z�/�4H��{�����/�e�%����x�	�0k�­%�"F�^��2}���C�H��RU��$���3A�l��x�P�*C�B����9P����6X(�6���חEȑ�3F�O����6ŷ�~���{���ҋ10�xh�����8$�qԏ@Tu�8��$.
�.�,k�G�����ϘM���?���zY��
�G=Rg�7���}F�"��ա��ts�,Tޓ)z�GsF8�V�FBӖ�*�)����4����4r� H��5�EqW�/f�%�۬�𛄓A��Eژ� Ă�� ¯�6����,oN"?����68N6�����wTn��%W_o=E���Փ�:��d�{�6�
'V�2^ �+�X!=Q�|h��L�X�=��u �&�,�3+
������6�r���a@ ����ePr�tp~��9�E��u�~�\�B�ϲU�W��.�(5���V�E0�a��,�*Ȕ�=�gW��y6���w3�?Ծ�Z�̏�c��"x|�ڝ=�M�5�ktr�W"���2W�R��|)LW�>�g��	ǄLgB���:q��%2-������e�Tԛhh?��F<BsZ�I��6��g���|,h�^��e�Eͽ�b������)o�=����և��?�>��H)�ct�I� ��ZD:��F��ZlL�.e�Ńݜ��G+���D�8���%�wrxԃV�3�Է���"K򡘣SH)�[:U|��L�P۪0y�2��� ���F�`.G.Xb>M����iy�sL�1�%�*������N	i�X LR	�}��F���J�>1�S(�ґE��:ij�Q�&��� L!�:�SF�nZ�x� 	�7(��$�P�J�y ��(���)h�q�ꉳ�;�x9T�m��
;ys��A6饄"�B�Tdu���,�lצ�	��xu��p���U� ���q�.�����D=Yԙ?�.����-@����$J\�̩���C�����
�z�K�чn->�� �Y�1������q�_|T�f%sS����Ư�s��iݻt
���j��A�P�O��(�|B-y8g�4�������C9@]F��}b�=n����l��O0��{i9�TT�d{z�D��	o0[x{?_FWz'�t-��o��Cj ֘�ҕ��n���+��$θ��w��p.�0�D��$����;u�<��􎿐-2Cw��7��_v �
A �H�aҥ�m>L�8�ٚG��8�pj��l"nK0٘�<���������ˏ�����ML�m������B��4Q�<6��ݸ :�i�:Y@��k(��X�Xꄪ����?��Sh�v/}��骞�LO=\9LrhP?���ҵ��-A����ʝK���{NgG�D�A�=�*��l�J�~n��e���txX����N8~�ȗ!�:�C�>�W.� ^�mR�v'��6U�`8��x����/�i�%�@����!yJ�r��(��e;H;�rn1Ů���ֆ���J�c"p�N������f�G����P��zd��������6�ݕ ��O�yv&��8~�ݱ-ne.ٿ�����S�92��.�?�S�B˹�-y�y�hY���t��U����������P2��^�Hiq����\Qi���0zi�+L5����:�Q�U!0��e���h��f`P^m
�L���GcA�����ug���V�������]�D6�v�e�ׯ�og���)Z(���{Sx*���V$?�~lk��!��a�3v!u��	�h�����N�H�K�ztM��?�[2$�dZod�+Y���.FZ-�`n�酸3���
��\;ߵ���ܢ���B��� �ƕ������P�Mb�6qA���T��y-qV��SU99�W�70�BL���L{f�g���4�O@�Ǌ �J�~�9&RG�6����gcc�B�A�[o�s#��R^ vN��r2`L<�G�u�*���%��u��.^c�(�	��[w /�E��x �II�6���w���i^�.��}��-�	,]	pD#��Պ�ҁ!���{q�%Ɗ�<����V�W��cB�&�@��@����d��] �(<uv��/��gt�/'Yi�M�,+��<;B]�Цa��'izS^M��;��5@t���j?x8���[�w\U���ju\L��������/�4��Ӡ���*@$�v��硊1P۱��M�%o��j���}uxqV�� ��	n�W=�:~�_?�zӝ�*��*�e���w��r�^L�R��Ӌ��xT+Z��u��j��ϣ�4��գt`���h�9��a�n�3�� ���&��Ǻ�̬�6����ݏ�ſ��ȕV��E��+Dڿ~^LsP�֍�%�`oAX�z��¬C��)_����2o6<�g�#��s��7Jr��!�Ew*Ck4x],�~������	?+��9be��er×'��,�F��E4���ݕ5�i�v�&r1^�[4�\�E�� #H����[ݩ��~�w�Pr��( �����3( ڽv!�\�O�`��1>�L�\h`>\~�.�9�ҊX���ʄ@Sc��ܯ��xa�O_p�-�H��?1?��a�z�5]-+f��2qh��'}��]�E;K{��J���Z�����N������n��1$���+��� �GDz��V�$�!�`�1%�Q�+]Z܋��V�$�ͬ�g��2�߰��q�G�6�5�,�ù������i)�=d�Y�����uԠ��K��B@B�KBDX��e�z����t��P���Jel5�� �����u���u��b|��e:����j�~��P�O�zXR�i�K���,:۝`��*�Z~cTp�s3 �ů"�)OI��C�XDs���`\|<
7-G)ٺa�o���	k�J�� �77iD5K�+���r��J�[�f���z+.A�JO���ULz�p�2�ǥ���3pu���d��8�4�}c���їO�>�6;1�$��b(�o+pY�-�cO�t���:<��X�d)� + ���(�4�d �}e�����%�"�m���؝��?C/���ZP"`�H)Ŋ��s�9}vD�7"���#AH������D������]�p=2��ޕz���ߨ� m��Db$�{���7zqMYm;_��]�t
'�D-P��2/H�4�,�ܜ����o/��t�Z=�m�{@��28�9��a���t���+t2"�]�1Ϛ�f(��e�Cr��:@�E�]FY±O"
�ro�փ����3!��>�U���_(5ǈG��ʣL��cc�
���Rʑfd��xN��ס6[���U��:�\����czM5�DS��?���r�f��������h���X����R��U�
?si����˰��F��{ל�ŬC�-�0f �R\��k�G�©��$.S{�}�g��F�x��B�c��j)����!2冥�Job�/y�gc�����`�e��Fe,��,�AE��3K
�Z-� r��<���ɶ�o�ѝ��yWEIς�z����)��R���4�x)L�H2t������JQ(��i�y�&~���&��/��$�����`�2DqA�u�v.ush~d�FƲ�8����X�Ŵ9+��p;А�*�@�E1cgYyrG_U��
�vM��]Յ?W�y	�A�b
�)��Q�U����̯��p�`\�N��#����>��<��<�ǉ~�<���x�M̚�qfu�п�%%����FB+]��[� PA����b�M����)"��H���#ԍ߻.��%6����J���&[T�V{]?�����	��ڈ4�t��OcA!�Lb�[M�j�E��v3g{a�u#�a���]#��/5	��P�1��c*�!�<�����Cy�XC?�s�#O��h����ƭ��#�Q�P<s�6b�*�*iz���ҍ�6�O��SX".��1EA$"o*%��V@��s���Kd�Y��&ο�7���	L��ˋ\��=]��y�eVI�+�&���ѫ{���s�rB�B%�����c�g�Mo��5B��22ߺ�'�+2j�n=�� �j�`Dߪ���넘#�}lg����١ I;�S*���4�;7�I�|�I���ɁkEPx8�`wK�s<{�j�K �W��\��)%G�2R���*�ޥ��Q�D��k�����9�D�i¼/�!j.)���U��o]� _��x�N�X��rBY�¹3�/m^{��mL�aZ��h%�� �*��<WR�4u������yL�q:�n��7�1�F��g�A�<��̳��5���׼<�عZ��N���'��������S���c	fАD1�ټ
ݭ<s�����)���t?D�Lsn�����A��$�F�@1����΋�����X�R,Z����FĊ�e��%�BC+�싅���<���cIy�$	�I����ב(���mRb6g�SG=�d���'�c^�8�aH��.����/�
ߍ�dK�|�����j� 4ĶnYv��{&�}�*R�ot����#`H�� �(�\��)�_��xJa�-W�w�P��eB�����B�	�q+Q��Ⅽ-h�m�
�n�mB�Z�)U��}@�Z<$��@��&s���%	��sy�!�����o����I2o��+�H���Y7~�ڸt�}��gS�c��'W(�z�g�څ�_F;�Ş�a�휏8��'��������U�*���M�\�Bo��eư��Y
��Z�^&6Kwݑ�9.	�Q���QS󦂢簌�^�����?��O᧲�sz}�V�n�u���K��6l�_3��p5U�7��v�7~5@[�$��s��1P��_"Y:��=���%�na�oKCJ�̅�}�Y�I!��<��
b���5,��m� �f����:O�������H26����Z|G��� Y
��j~��&U�!�+t�4�����R|����Ͱ���W]�^^��1��Ut��,+�-�S��ɆS�b���n
P!c8�����qN;���f�~�z�"r�(Q�~��,0.��*��V�F���]���E	7�r�������&�CBq�~�`	�17\Tg��o(0��~Rj��C�]]���S��G��C�]�ܭ�^4�cc��{D��Aj��k��������vU�y���4�WKۍE4�A��X�ND�l��N�`d',n	/
ə��|z�E,�W×|Ɗvg�x�o�Q�HScKn7h�T��]J��c��73���:�m��\gc=9a'��Ђ騡L墡5���-2M�$�6�9���n�\��[Y|	6PB��0�˱�����(L�4�3lP�
�|^��}�
B�ս���a�.UpI��r,�����yŪ��p]ʝ�CCS�xvw��A�=(%���E������<�T s=u!��P6^����B��O٫t�@���Ι�"�(�e$q�x1*�3/&�(�v�T��k�����i'��>�UY5��@O�#��,c�Xr^�����{�����!	��No���n�0)�w*��R�h�u�O����:���s��I�2�o�������Ѯ�R��[�'�|�}�љ;޺�ޫv���w��D������Gt����:��_�o	S��c�U��>dݺtI��Tw	W���$t�!%rYc��<�k!Umu� ���O�T �����[�����O@*�W!�R�X����ɡ5���j���8w�>P�a��E��ۼ�FC�u?�,A��Ɗ����')�")9h�Zw+,���""�=��L����5e����ٸ"�s��`�%������{4���k˜�`m���c������&�7��s��Rv��.���]̖U��A~�Rz�O7�w�l�˵�4b��p�Y�	���V�;���蜐����?�R0��\Dp �1y��܄���ʯK�C�����6S0��3D�j\JM�0��%c�BU(OH��;�??2�J�!�4�d6TGjټS���68�M�!x˧����oD�BE�Q53[Q���q�MVh�1}&a8۸w��Y 	�`_�lڦ�H�m8!v��\��k��Ryf����A�����#����'��f������/��F�za�?'�	i����*�.;�mL�ĳ���]>��64�=��;�&��
y�������rT8�Q�y�jAʳi�mؕQL�����p��<��15 ���pO�����bG/Ԓ���ڪ�_S��ڨ���>��,u�{�Aj�w֟S2عj�	�&���ys�����ƃ�Q��=g��c��d]9>���/3�5~��᤻��
C�&��>4ϩ������e������;VM���RNT���yvE`;��4��3�K�s/4��{�%�#
�f�|�>���d�F?NA_�Gc)
0]���~i��B񭳣 ��P�-���-���Fk*i�B�!h>��"��R�ك��w�}^{���gϳa�p�c�� �7
���R(�;�O�n�F��Q-�q,�#��B��2W�w�L�7�|c�B���|0���ڦ�����"�$5~༟�cq aP�<�1�m+H�5r��Ӿ�H�OT���b��٘��.w���׻%�hR��?}T1��ה`���s�?�����K��A���x7�X���'z��b8O�n���<�}&�`��s�G�;���_���w|#zx��P�%�֦���ٜ�+�s_#٥�`:�"�ڸ���%�O�_�'0��ƺ}t����^2mY����`�y����
���>�_\	Ӧt�&wm��Ν��Q�����n��F�lА7w�Q#v&���y�V��qGO����J�!5�m��*<w2ؒ��i|$<�n�cP��j�}z\���ʹ��I#�Sӫ�V���_T''��'�?������|숴9q�N�p�����<���ڀ���L@����hh=ng�˙�^+�	���%��?�6M������c��dإ��5~Q�yI�{�[�l|&�S�4K�#��\�G'��AuV����a�M�9�g���Ss���ꅝ��+f꟱.�=��4�O \P5��
"�8�ײ]ϕ�XS����#J��$���xw�aHWF'�hp61w��"��*,�p�^ [��0��Q�̀��`c���iڭHe�\&%g	����p�
�`$fF����q�*�-�F(#@h�|�rG(k����sX~� �=j7(�aRK�������$ �;S�s+|p�1�\�W�	��'
���^,l�t��ugy:�I?>��Zs_�)E%/
���١L��O��A�8{�
�XR�=T�5�u��`�j)�NW"M�.{9��+���eL�O�0�ϝ)U1S�'��|��~r�-x݊�#J?Akv�h�_�P_i��c�x���S��9"Ur?Fҡ��ch���`������;��l(��{^kcP*J�K��ْܾ�P��óF0�ab6�+��j�6���$���8�qz����Aq����O���k�M��XaE�x�b?5��
�g�\Xi����I�nx��Q����@6��utj[����ݜ1� *�-R�����g�:���q�c�m�5C�=d=s#R�Rߐ	����>)Mz�MW�R%�l�Y	����t����� ��04HΦ]�e�OM��!�s���?3z\!��ZaWxge-��]�f
I�����������t5
��7#it�~.2S�n�\a��z�;�!7�^��O�.�Z���lg��J��xŜ��\{�0T��7���M��YA�Uס%���݌E��ގ�H�΀��Dv�������B��	2h�+���3�/xB2�B���5 0I�\4�w��'YI�veZy_�.�)�� !,LB+��N!���Cګk�efKy������2'���܏�R����{�xp��~@PhU*���?����V �	҅wr9�1�ƱJ2)Tsӯ9�R�gހ�G�V��Cl	��kź�?� \k]9w�ϯ��C� ��:;aŹoX�@��"���]�1C�K�T��r���]�b��<�:M�������j~[41�a]�ߦ��/ϭ����3��Xw�
��8���,��E�p]MQL3Ѣ�3����G���'T��$D労 )�u��F�e�@ϋ�{����z��_ �et�"cp������дiHU:�I���Gi甐��頿�=���=+H-'(˞�N�ں�b�����<�#��F�,Veٗ\�nu�U�X��LK��^Z���
V�xa�JX�	�N|.� нI �������p~�?T���B݋����둯��D������B��<k_T"�s�rm��M���؅�E�ՙ��x�f�e�!i(�C�B6Ը��2�`����m�:��b`S"�;"�)��ۍ� ~w��{�1��,�rW�qXc��ࠎ�RGT��)ab� ��H����Y�X�X-<�O��Oo�C�;_ř�q�B�`<_�H��a4S�e [��h�9��'��5,hN����^1�b`X��2
r��P���H��(���QBw3�uK���6&�iu({��`c�������vI)���0�6!�ܢ��?z�n�7Iz������	u��`�O"	�d�J�&K����vi�/���C=� 
I�6�)v>L��t�1J�8���y`���ۇo��\I�#��}��a�v�)�O�SC�Ʉ��J��jL">&	�
����:W���A!}��t��r%�@nj�j��v�y�5����-b����V�٢��t|e.E�Y���Z���֭�Ii:?���論� =�}Ok��Ri��xf�. Q$Z�����pzt ����`��C�0yI͔@l���!<�I��"ް�����4fٔܿ/�,;�������S���p����&��Ȩ�8Avu�� �nȗ�N̬�V�0c;GJ[*[!�I�	D6��^ྲ�3�0u�$��)\��%����O��J�r>���Ù����\w�jQ�[l�2'�z̕`�H���4�"��N�*5L��G�8��ֳ��	�H�0	"�,�^��39-o��iE�ٲX�E��
�/JQ�����'���Sb�`ni�â�Š[~9�J~Oz�<W/�pN���4��sH�}n�&�/1�0�
NC��Yf�8@*u�r�jAp��=��%�<�0�f�� M�::z�G�\�
[�|~��|�̍F8=���,,¬ʍ̧�I�J���
ҹ�mM �(Aq�Syf��;-�[��@��h�|[n�X���n:���*�^�{����iڜzh�DR��^�?�X�H�.�aDO���褿
D���H~8@̮�ķgb0��GRv��d�r��!�{8�a�x��w�[�"V����XL�6��>���E�b�:Tl�-_����QıX[�b�$t�"�M ����xG�w8�vIjۯ����44�n<e�x�Z�Q���8s����.�>�ܓ��6�w�.H���f:�Ր0�������&�G-�a!��|Wϫh�lC-)1b��b|�	3$@��%�*�с��!Y�%�M)R}�����y�Aޢ׈m�z0�DA��,-k!(]��¢�9)���{q�0V&����#G�_Պ�b��������Q]��t�N|O	���6�'7 3B)\
s�w~�H/�+�Yt=�/�]�4����N=Ք���߭K,�8�]8?�?�*������0�N�F���A����(*��<�q�#_�9?�9�7��2I��Q�o ��Ia�[���7�Bg(e<��F�y6Nv,���>��XS�o�eь]�?��U&�w����T⊢��Vk/���Zl�O(�DD9o��K��=:��k{C�I��&x�����wOM-d'�Tҟ��0��[c*z�0 �n�T�X��l3)9�;�����5'��X�'Υ�[�ӳ�,)DV�����]>�H�&��������%�[��J��5����ހ���L��7mK"Ss�燆Ԅ6yþ-��de$����!;x��eA"j���`=���
��l�c	����(�ZbL��ߓ��p����mʌ� =�Q�д�]g��Q���S������G��,����л{) ���&7�5��Rw�%�gd8��� ^��1�k��b�	���<�T$�>�D�`�9��}���vZk�*�#l�!/RvW�"@Ƃ3#��
�q|Jw��㪨���X�)���-X�	3	��h�eY�R#I4.���;O������N��IӺ6��!1Wcѳ%�S�'�iCb�q�Vf�YZzب���׬���ߠ�j�h�N��y�ݶ�@��D#��;K�eo+%�SŅ%�u1��h��R*q�ZM�?��j=��׎Y)V
�����s�RP�3"}&xh�����it��.,�>������j3@!k�C��rc�ac��N%:�_����h�6�ET���e��b����~ܲ~��]BX���PN�@�%�M.���ԩ���]
��1�~��&$�!;u�4,�B��lғ��O�>�>�	�Ի�L�z�Q:q$�����S7�'�5;��)����缑k�],�] 2m���v���Zɘ}1�o������!<.��0�h�uo/'�+�w%݈#h͡�����j�0�O�D��:#�翵G��`���y��o�����hte UC�טhb��Ѩ1�R-Vm	Q��MO���ȃu%��(�z]�!I~+���44���a�3p�n��T�kO&���Sz�+�����.��!I�L��֌\]�t9rު�@x��7�\t��#ЛM!������v��d����Q%"�~�N,��� �ߢ�_��~K�����7o�:WA��p&`�pnl����ѡd&��Kh�Wצ��"#�S�t 5c��`�����7�.�h�ڣڟ�<�1�#]`,��h����~�m1�n;�W�}��Bӗ��d�P[l�pZ�/��˴:�f�a'I�\�x�>�� ���gM��L-��y�#�!��D��+i7��E�|.i�"�)��l����l>�f���XXY_����j[�Lm�$�l	˦Y�6 ����G�J�:q���2�����{T���Ggf5�$$~�|�X��zw���l9S�T�l��#!6�s��)�����q������?sf�B}\�[e}(��7v� �p<� ����9Lź�!Έ��ؽc�`Z��>]�s3s�3=�X���*��H\�[�Ļ�R��+ͮ���v"�����/8	����-	���1M���-�f��.<�W�S��I�c���hwA�k�<��ֲ�>W��m ����}�w��Y!(�<��������3P"��������b]_`��D-��(-0ܒ8 ��Q�b��Yc���P��&�G�[��3j���It�G^G�CĎ�`�v��qn4˫�)����9d�r�c
p�Љ��#��G�5����ϔ틃v'�ħRs�O�����~kE���wii����=O80�.O�=�H巺y��di�q	��x}�Ő��&�2W�i��x�lK�y�`;���F��o���]�����G��{;��r� �Mx[�>�ge�
�	�3�8�}�v��L�dF]����t��ٌ���h7޿L�Aɵ� R��؍�^���H�);�y|�_�O��{'�I������Φ{	:_���##h�k��
z+�f�f�^{�)��ìA�	#����Ϭ˨����l�)s*���¹Yz꣒O`x��{ ]����i�>��3L0@��~�
����1t����b�?"��~2oX~�wq��z+�`cO��܅��]u{]��|��|��Ѽ��`k����ۊ|����7�Y�$h�'�f%jN��Iu�����@��$]�z�"*wzg����yF�@�����|ƩV�x�y=�5� ���	��M�F1�4p�"}�="���cٵ�:�%o���1�1���V�?S:B���Ж�-���]\�˳�S�S(�^�,Q�A��q2����3h
>n�<AB?s-*w+�Q�%)�J x�^�"�n]`�x�N�Dބ\��-�i��-�� �\�9�PH}�;ah7����{�w��=��n�M
�G�\���G�a�_㪲���z��t�{�XR�����滼����{�����YŞ�� ��}3?h&Bj�,��@݉�m �XR:�xL;�
%�G�wQ� o�;ܓݠ��e��m
�t��ǿiW��QR���-X���ɑIC��Z���X��U�ຝ@�ֵ�9����jm���C�K�H��X!�Γ�٤Q,M�(�`���T�ʒ��(�U�@R`�J�ͻB�SO6NZ#V�����b�u�T(Z0�(�fڋÿ��BF��nD�ޥ(n�e��-�/����г�f��ȧ�ȗp:kP�5L%z�ϣ.��3���eak�Sj}x�k�\ɖ����rZl(��L�؇��K��X��eYB�1�Am	��`����ߓL(��d�V7�뀍�����N����5�ʳ���>��:���C�	)�r�L� [q5�l�J�f{Ϭ~r�c���ǐ7�%�|�rB30��i �N���ҩ��ڄx�*��=*?��g��=)�[" x��8��otsU��WP�K~0[��e��l�k�|z�=N��ʮ����H`n�����RE�3}vԅ>�ڟӸ��x��@&��b��bzca�#��慤�:�{1�U�4:@�a���s'6_��l���tE����>��U���'��z�uʁ�N�"�q^��?{Qν��'KP�Q�ƞ��I��uN�{�a?>�~>����|�P��xf�T�+����f�\m&�[g/AY,q1�P���{�h>;����8�fĎB]R�r���ۊ�4"k��hNh+?٘���2����-��1��
�M���w�j4
{ F��%s�g8��9�RtZҹ�p`�Cx���F}�����O�V@�}��%b #�􍎣��}���۟K�V���cL͞�
6&�zCL��G�p�%HH���*��av���9���Y�-@@�3=�?%��L��f����� ����50���� �'z�ρ�\�f�Pu�
i�y,ׄ�@\r�yb�K|�ox�3��w��+R`�G/z E�B��GWQXΡ���x�{wK�ƱTu��je��]3�3?��B��I�I�V�Q���;@�Դ���Y����N�k��X��Uv������j��jb��1Rh���b8$������ǩ�s�ШH�*�hK�\	N��[2nְ���������ak����bK�1~ܚ���/�F����[��I�	�ǚsfɣo<hCa	�iJ	fSK#��� �*���%���c��iԡ:�|k�RDO��]��}���߫���=�����2=Z�mN���� ��}����'ظ���_�{�>�L��*$�"J?���v����B�$O'ӛB�P#�[�M[�n�Mw�0v%m�8���9}*8��/�Ds�p�(��q߱w`��Z��0o � Xn�Ɵ�e̺P1n$���S�婠F�G'�VK"G�tg���n�3r(�?�.���
�}G�Wr$�
S���=�+�bj�t<'<\���� ��7�C�T�+GV�QfW�����Ê'�Q,�O�TȬc�ݞx�#���!��5;���C�h���m��7oP�g�Nw�ҥ6�|�"�� ˳s�ӷ���a�t�!o����4�R���B�t������嬊����Qͬ"�|%v*�x��pG��갪�UD}c�89?�g�P�;`��T!*��d�p��/bCr�+����[��Q5�[���ژ�� � �������0�M[�C91"��(es�o�^� �@[���p���E ��<����w@�E~��x�1�K�퐦�B�wg��Tf���]��h�c��^�� rx��,�;��ѓaT�����
B��IL�i����XA?����Q*~�v��:oH1]E� ��_�'�B�	�;��jN>١M�l�}E�,گ����W�3�6�lQ�b8���X�Ъ�Q"�p���v��j�aP{�վ^AB^�����h)&�z����3_@�x�Pd�|��a��;{z��<8�+���C�	�K&��X�s-yqʏ	��j
z�������aq����5�?�`���V��]��E�>��d�BV��.Ed����g���cI��{WO��}D�{`�$M��X��}HSD�<n:���l@1�5����c�^/�j�xsgA���	�#	���y��Iz���>?�X�L(�3�/�L�em�E�r��@w�ے�ڽ����2��Lse]Ϋy��`��,"���� Q(�q������J������?tް�N*(e��!*�ug�����Y��)Wk~���n�*�,�-%W�gJn����-��ySZS��_G���I7��I�6�A���Y��uV�$H���Ɛ���v_CMqg}Z8,�"ń�
��B!g�zī�&�j)�z���|�<v��.yB��^	���JV���i-�
��󩐀��iz�8@v�(����;��t8t�o�J;�$._.�_Q�� ��iGy��=<�*�a���j:TL��'�W�Z
(&��>0�3�z\�_��Epg��k-A;�|���&�iY�X[��,����D����߆A����W����|¬y��gMXJॣ��|�����,y���E#	�Ϫ3�İ���zUZ�&�#�F�& 	ծ�kO�;��V��2�t/�u����mx���I�+�r��-�1�����Q�l��{$(gu�}������
{`M@�xmݜ� l�?j�*������1/c)�y��d� �4����M ����K� ��c��d٨)���kUxJ�6mN�W�#�&z�Ш�>mL��J������JRD��Q�FG�C��_�̥�bfIVc���\�+��-%kH���X��F������C)WrR���+����ď�
�s��˻�,gr�� s�<���T*�9�ߋ(�� �nZ}N%�o��ڱ���֢��?��|p�Q�;�N�P;�\:��m�a�꽂���L�C��޳����F2.��U��X���M����i�,Me��x�y�;&������7j#����|����S�2��_Z�u�!=&	��m�&[j�E��-IgB0+jI�U肛*?��:��ט&�!/���R�f�g[N�D�=�������[��m%��l��5T���-y�e��Dp��۠o���uSJ���nɋU�ǫ�$�4^�h��2<S7���{�E�L� L9j�do��h4�+_�m�$�ko%eh�K[կH�`���e�i�������+�x�1���m�,��r�#
dsN��b�-Ѻ�f�_?�P�f���=D��%۸ӫ���5�D|)Y��M~���Xn��kq�Wd
R�+O\m�� �	���[2��"�=��oJ��%II<�dVˆ"��tTx�T*@g�#*q��iṆ�8w�k}]k��k^��b �!a�^uڢ{y��$��H0�}*����Y;g��0��/�rؘ:I2?;�鯯`��n��s(�n%:��Xȁ��|��l<:A�v����V�`���4�oP�ϊ�oѨ-������'c�=ɐ�8!���	3U_N��p�*G�/�9;:JO�*����>�R����(�"Z�0�q�2�=����b~7�;�@�>)e����1Cd��G�lu��IpN��9�k�o*��d9{����ע;��@��-g���&�u�4]�8g��ݱ�tI:���ȘW�^�y��m�v��W�����U���gU��ќX2�+�b�G�mʺ�^�_�`��88Y-��r�y��f��Hd �>�N}�(c'8���tg��qaynr�(;Lo�q�?	N��I�h��n�K�[�K�����������$���Ie��N�O��(N��q�e'1�S�^�v��K8����fm�K
 �,������w&�����j���+=|W�ש��M>_.���<C1 ���^vO�B��������aJ���@OKj�9!� _a-rfԙ2e���:z�5��Ί��^2�!^J�\�2���A�k(��Lů������:*F��xw�Q��+Ũ��9�b$�-�d>�!l���lQr��|&�c�N��=����������.�����ho�\���B�y���S�Գ\{z�#��JG+��%L�k��yW*S� ��q^X��Ww�����mM�|�Mq�	�W��(�S#���2�n��ą��ZU���f���:Əh��{�|Y�lO�iA�1C!��l���S��y�R�j����yxCs4g�f|�@��"Ϩhξp�� 3&��N-{i�	(�>`)��\��A�!R��A���~w��T�	G�(�� )�-y�,�9��,*U�{�r�mPDM -'�^,���!�k���_��au��d�Y,�J��gY�n�z"�C-�p5�¤�D�/9�u�ò�r+���f���ቪ)�p�t�Dÿ�NZ550��EO�4�?m�5D�hu�4��>rv�j��M&Y��T���d:W���A�3���	��%�Deg���(���������E���%��.��X:�%�i1�m��V�@��l?AO�1x��#�9�x���/�mXR���548g3��;ԁ�Vg��Ϯ��k��cc���َ�ݜ�"!L��𯎺 ����.�[��2�9��o��X�no��n����o����v->]D@rA5Kg�aKoY�Aј�U�yn���ڱr:�e�zGܦE��B$q�*l������_��Uv�qLd�y�r��a6s� b`�"��zJEʸr�U+)�{_�a�H`3�pf�X��4?XX�5Q�(Ug۠�K���l�Q�^� �~���4K��ԋ�l��S?���Q\6� �Q1�U$������| ��Zr�`]i��~�!�ڇ1G궉v����J�?9~�z�X�5��R@ܝ����8S]����T.�����?p�]�RbY�tY'V����C�S�<�s��y�=��|���Hm���{��{�R{2�v�=ϰ��6_��N<�s��o�	_�gM�W�EB�^>cf�����P]!6�n�9�[6�3�[;C^'�*I�P�+�F㐅en����J�/���Ŗ�96���2
M�/[@�3��u��
�]jt��֘�w�b����1]�	�^g��mn���X�L��WTi:����n4��"j���$ƅ����[�ʀY$�>4�Ɯ�Y�:�sΫ[Q��J�ww�,�����F�H�?L��$�A�����4��J���T�ճ����h[����@����Z	x_���}����Q�uH:U�
��k�=ڙ����f3�#x��g�*R��,��PSJڪ����	�T�Q{�v;6=I� ���ȼ�FAu�ǃy7��T���x�L���5��o��������
:Q�4b;yғ?"
����@; �5!��j;.n���K�Q�� ��,�cۣ�����KO�`���,z����(!{U)�c�ɜl-6��M�3g3��3H'�S��_��9]��Y?������u� �k�� \8��MԃmY��Yo'�`�*� ��{'���	Ug��z�D����������P��+���f+F��.��ͱ�	{	ڸg�=oI?�}a	���7��dJ�(��r=�c��t��>�z�^�6�u���Zʠ��5���!DF�N��`�(w�,%R����Ej�3�s��+ӛ\ʷ�e5~{Hǿ�;לXd��H<
;`)�d��@���z!�7���TJ�Q�Zi9�9���b\��GLWp���cܱ�Ь�湚q]72��0��<�������E��"P��"y��a���BH.]����5p:���؉��Ƭ�8�s�l���5H|�)}f��?�[y��^���֓-C᥅���a�퉅���`�34`���-���7����˃��vD�@�M���ΕV�{�y�W6��+�]*�g6~�h$&[˰4�Y�@�%!ƥ×�?�̡J�F!SOoK��_5�	q�6�&;r;����1�h� 7�ecj)�*W�ޏ���*ш�؃�A�h��>'m}��<����ʒ���~���!a��Hr��9I�fS�	�S!���j.�pMkY#��^6�ts�L񎜰�n è����E�j� =G�O�e��S2��F�ô �m�ʥ@T%e_���c7�:�Ǉ�Κ�A��!+d�u�?`<+@1]��rb1��Վ}ˑ�M�	�:��#1=�.φ�N��8Cp��q)T2���|Zr���P�A^z��m�Y�x���x��'�'[ׁ<(�q�+B�1����=Y�~BB��`zOC-I�}�G�;��p!A$��1n��e�=3(����f�TE^T��}Pe�L9qP�;�g����_��|c#^�]飐�e����>ʔm����u��dG������P���^��?���r� �*���F��A��|s΍2�� ]6�a��l�Ȇta6��!���vj�����W�� �b�H���������NPq�l�"�h9��o���^�/!� t��aLt�2l����ibY�9n�]@pZX�=�o�Q^dZ�e��3��j���қx�������,�U@J̚dr! i�~������t�50U%��!;h���tw����C���ZY6����^b���0<=�?_��O��}��k�vhZ3���^<1ihX���AFB�������kM�V�>�4�����Sɦy铯�Ė��$���o)�_����u��H������	��h5��P�����9h���Hx�	{tșWHC��m*v����r2\�|�e��%{��K�
�Y�,� `��9�V�x[ e�&�� �C`�fЇ賫��%�9��
�ӗr�qc�̏��Mg���H�]���X"��U�ϾD��;8��{Jf�=+YZO�c�s�����G�2�D��K� �/D6��ڰP�H<�y'����%�g_�'����\y��h�r��1ׇ��9d�Q"�k��0�I�e3�۝�)<����6P�ϥ�Q���L���!J,Yo��-�
49�Y��������xϾ^�v�}��3O�:�f�f�A�#���|���bТo�'r"؀<�ml��|�Ir�cF���pz��L��p�i�D��	��H�X�+<U�[W͹(�����.�(Rbڂ�"�"�c-��dD8�S"fGA�0����=�k�,y�}:^�J�+��nbZ>7i�h��(8�m�ޭ����6�b�����U��n��|�����sTJ��g[^��o�}�Cg�Fې�Rי�A�r��Kl�o��E����Q)�U����1�d����7���,�3yw�9?Nmy�#l�f�t���MR�� ������E�Т�ع�"#��c֗��2�N����V$q��+�������܂�f4�X<���`-�~/���-�w��M? �1��
���LM�g$@�U�YKE�<Qc&J	}�$� ���<|p,�j�?W[B(���۩��>.��s��.�j�奈��&�<�w\m8��S��<�5�aK����������N,�+A[�q��By�0ME��2YG��b�1��<C�!ֵ r1�3�F���ma[�!�Y̡&�[��p��謁)��7lz���#r�D���gk=��A�A��3�YE�hгl�c!m��I�������/�����IoQb�e]��i����V[(DwMo�V+��V��ln�	f��H��Td���}�^km#�;�=�_���Sb�%O>�O�TT8���7`�^
�A5�N&�%p�M�CM ����۳�˃�"���ܥe�G|�}���F{���]�2y��2���OJ��(�c.��<�-��J EJ�O!IFÅ�'A"(���RY֞�t=�
�%�~rl�.��(-`�_޲��A�0+�.��5�o3|�Ӈ&R����%!	�gZ�������("���^7�t�,(��V{jZu�˩���LB��a�����2Ю�|��K:�G҃ӵM�������3Ia{���G�{k³�(��S�A=���wW��bx�&�3�^����W L.�WL���V�����J{���?ǫ�N�<t9�����6~�O�f�g�VH4�FHB��r�t���ٷ�췽��'�KW�I/���B�I]��\eM��r�������)��LZ�����E���ktңC�M�;b����m8͈zʇ4}�FO
;r���R��@8�u��('0m�0�x�ʂ[��޾��Tru(yjCɡ�5�W�UBQ=lK��`��G��t5	�iE�Z1k�����PZف5X<A��� ,�'��=%�D&����V~~<�+g"8xx�׺�*N�R���7(�����d��s{��GØxn�h��y��O�+��/���F&���/�q��0V�
pK����]���?�(�4%�Nͫ���NUM�����d���T�[�.��]�t�ZÆTp�^!Ҩ,[(��I32�y��$�"蓱��~�%�����U$��1y�j�fL�S?JAn���NV����4��U��S��? ��� �WrlLd�����-C{�ˍ�=��<�ſߞ\����/��l4jӡ8K�%������W�'�j#١^�i��S�P�0���u6�N����1�o�y�DT�_�Q�\F_�;��@�H1�2vR�����eܲɴ1�0���/�E%�+0b�vL?]���,֛�)8�$�*����Ж�6!�]���]�/xn�u?���ݶY�n�Of�1ۭU`z����+�L���ۥ1}IDD���RU��]��AHm6�NaJMwA�mLϭ����! ��^��p���l"��T�vmL�I4�4ӊj�l�S�8�%�a��{������_ƃ��_�ڦ��/+�+7��
��딘�Z؞p��\J���@{����I���PK�[Y��@�f&�١8_��Ifi6-z4�N�k||����ퟷ��A� ���pB���u@�d�����܈8s����VTui-��SG` ��n�y(�؁B_�:~l�ņ�is��'2��q���i�;Y�~�\)zޤ�X��/^�Lh�����~�0�Gሶ�e�ɹp���B���A��9�AA�(�Us��u2�ԁ>���ϖb`�2;�0��-@KS7����Q���A�%B�Mg��\W�%�L9�9;�qV�%d���P�4oK~ߕ�"Ւz�IO��Y0�V	���1�� ��I#觪IB7���E����=� ��L��-��%8�:\����m�y4�^>��H���vy��q�9���|1g�uE��_+�|�D���7Z�e�x94|g�6O����"g�1~X��7j&�R�s�F�-���t)�+��e0tn�W�����*/BT���YV1��4��$�+�V剩Jw��e�j�����"� ;���G��w���4V����}�	}A�J;�.��SI����!�\箷0|/����F���-�ہ�D��W��}����Ϋ*�n���/��<�_��D��?�Yvլ��X�����*c�q�Mj��/A .�c`�������_<{�������蹡�A��5낇��_b v�3��%��N\��.�g�5
%Fo��RQ����=�SQ"~~Z���Zכ!� ����h7�:�Ł�%��q��p�l:)��7��5�9�ʿس*n�ZZ17�^&�0��=n��_cf�z�P\1�ݛ+���A������ޥ����/6�*���+H�J��ᐚ�	�X�[�;�����-�6D#��E�殒.�r��<Y���bv*�����S$�IR/p_s�7�>���٠P�H+��=����[`Āc�>FM�ڮw~���#
 l�b�6�@�%�@�x��t�Y�Jl�5K9/'l<���������^�9�^3��Qx
�>���O&5�j�UĿGoZ��6 �P=�Hl!/�1D����,�֬���ݙClT��� -&e͂ȅ��g�!��)T7���U���^m�O���~ξg�L2��ш�]-f��r��"h��T���&��e_KQ�6wI���]*�v��`pNɺ�Yٯ%CU0A�� �#��Ç�1"���/���0E���jՀ��cuO@��t|����9G@�S�[ߦ�2�v=:�j�H���f�սH	E�%����~+z���.�@�U�!���+����x�H��
��#`#.��e
�Y t�MF���U�4����E?��h)��s�"7g�ub� �xe-��*�<i�As+Y��@ҍ��'[00�qs���z���;,��?�@3��5�u����`��:��Ϛ�n5ĭxOB暊0c���@ч�N�/��(Wy�X��j�q��!��(:��A����qT;D�`wU;�X1pߚ�~�ͼ�|o1Q��L�~������i���㐸=�%7Zܗ�Ǵ������O��n�D�T Z��/����@�99YQ.�r�7�T�Q5T/��<����6�� �Q���(�|��d�}B�&��/q�l��h2������zSQmIP2+Ú�Z�T��ʵV$;1Mo٥��<���覃�&>DπAp��J��
����#{�V��t��kQJJ��mG�)Q5V?��[xІ�r��CJ�c�o�?N�Ψ:�,�9��6�I/��f��k���0���gG`�xCȽ^�C��#��9�#�aӌ��d�A" �B��S�H�6
<q��$J��V_E�#��(��u|�	�njd�i4h«��n@�R>Bf�3L�*N��������]IE7 +4Q	T$�E�S�2�a�{Db�W�ޚ4�>wGJB+4li�4�������+;��2p~���l���䦇%��w�&��m`1bA��.��0ť -0�.���;����S����]4r[O����k�n'c2��4VSK��������7�V��A��X��2�8��7��8@෠� W�Kx�����rm����Y�`P��x�3<kG&HY;��d�O��{�Yv�K0���cs����b�i3S�(�.��4������wy��ww�SC���Y�a}�e�GHE{]�������軭u�T �`y��*3�S.���-�m#
4�	�M�����&!�A�X?x\I�V��g���Ke�p�Kqԭߤ|�{�����r*ut5G�������)I��k�I�	wh9�q6Ad8#xL4�X�x�B�2\i2����`?#�TZ��v4 t9�H��7��y�>{�04X��J%��Z�b+���Ϛ�_��G��h��m{�u��jDUI7(�n�R��ߗx�eD6g_Y?M&��z5忂S?�d�l��PO�X���������ܻx� ş6X�2�.?��A��� #~���4j�M@��i�������L�\��6!����o�p�}l�h�\�����m������M�����j( �9��#����G�Q�
���D݃�@2�j2���_�d�Kօt�Z|�̦�����)�VD*d�Z�t�$Ͻ�e�������0��޺�� (��!�'g�ʕ0�&�xS�R
��l1*g�V���>YB��Ө���J��Oe.>��#���8��(I���b��o�w��Xǽ�s���A��+3F����yn�pQul g9�//���%jo!�it(���4��`�i�Z��i{dN����(�T�:<��@��-t�r�^?�vd�	�d-�^�-�;g��}���OO©K���:�E��T�_���3�rޫx������pk-/]�iw��Β�~_�҅����S�������6���z>��z&9EǓ�v��n�¯~�?*��4��3�Ig�[���_�׃�8��@��'��(B|�T];[��yZ0�GyHW���2�X���[��>"�v6&U�jJ�%3m����^�pr��S��,5�3��ʟݔV)��Ho7ʐ���׵Ю�ar���f�D\=�vb��`�,[S�
��:߾�n_#_t;�(L�-� �z�T~޲5���
R�z��y�JBj�`m�����q���i�ԇ�	1E
�����*���A�O������=&`B��V9V{-Z�1`/L���(��vQwN�-L�'1qc���N?����WV���nu�7���4�ߕ������cݰ�D�{t�:ˏ9�*��~�G����h0B�s~?`s��]��Zn%�TI�!�4�"��b�����Ra;K����'re��ߺ&%��U粎�J��A3�њK�W� +��з���\#ށ[�VC�R���_(��o Be2y2^xV6g�Y�u<���2�z%s�'"%�=K�}�،�!Y�����c'J���^�j�R]!��}�*�L��2����7�8ps�~a:r���_�c\+z���^-�>��ꦬ�J�z�Nv��3sI��$C����h��x��%yt��~-�8�>��[m)�nS�jcn+��=>����v�&�p�M
��*w�>���M�_���*�2t���d�����Wg�5�Q�S�����i�U5iD��,�}�,�nm�oG��<�@@�Ҭ:c�f��U/$��72{�X�J�-F�tX��Y�1%o��2cZ$�v�GԠ�-�wùH6%��u�h��̒*e�/��Zʷ�N�UP������\ 9w�C0
0!�ν�R��]i��J�b��R�ڍ�����n��+`'1�����d�5_���X��˙oYp����(�7�վY�?<�����]��͘�e������\�򹦺����s��ܦ$f|�}�Dn�t��+��YM�۟k���_��8���!��0��D����}p/�#����� ���2���aa?��TV�NW��~��c����j�1�����k���,��sW���N���o��G z���~)�bP�E]�=$��4��^n
/W�',P��w�'D�p�"��u��[̓�	7��(R��G�����c�t��A�hc}1H��ҝ��$�ig��ǎ��+:	 f^G/��_��������	I�[��e��k�|/���gٰL�;/��jo^�n�l)47��Ł�n�Ƿj�Y���^c�U�Cղa;4�!8h8�s,�M���|�������Ӫ\�D�SK�oP�=���^�ȟq"Q��[ȜlY�#ěp���P�}Q�����e��r�rX��L*%;3a�_�O�f7L `�n�Qv t����j����&n۱������}�p:1mB��S���`Y&.��gΕ��&3�3Y�W�1��� $����P$�y��*�+n�>?�������$��N/�:/-ӱ��e���
���rn8�w��g%T0�VC�+��nX6����^�m2vb�H�Ԛ���EoP���/$V+%�~,wu;o3� �Aw�R� ��sڵ�翷[�.�v����<]�]|��L��X���ɥ�ާ�8��qGƵ��9�`���5aq_0���h*}�h�ʢC�
�Wn�;���4Fw�g���`򎼯���WTM~yK{�b!���U2�n�ty�|uZ����HQ/a��Pp����&��g�=��q�oY�	jQ�Vb���S�M��.�$JF����X�Rsn� 1�����]�zذ��2N�#����P�CD�¨�Y� ɉ�ʌ�"�9]N
�t��x�~�����_����¤���I
���EN����;��xO%뻺͒����@l��DW��������5S�m����0M->����ꊮ|y<�]$P����R7�p�WP��G+{����ځ����)���4r��|��9�� �M�S�;��6r�)�JC�k���:}�����/��!�csup`��ت�B���+�t��[~��n:�O�	��h�V$��Ԃ��7�y���-
}0��֌.�mw�A���ky,e��U7ݱ&oF9q�a��xUe�GT��E#��j��A��D�_ّ�=���뚠��j����pI����UU��D���v1�
��@f ����Xg^gR��+�[�t�J�8�!|�-�~��s#_u����w�tnP�HA�lT�%-���E����JF}�+hL,@���=�y6���P���
����q_>�����n�f�*�y�#l��K�jF,A�1泰��K�ȖZ}�G�0 � d�uW���cUϴq��58�ڲ�7H��F��=�E	�~��2��I����īx��d�sܒ=LU� W�a�ب3e�r�>pŊ#��F�iyB��Q����6���O�'�@Y�YϚ+�,!�mbB�,��o5V���{�Oɜ�s)��7�]�熩����,d#�j�Xb �㎉�Y-����f�a/U���=�
%�Z���5���2���Zb�V���oQ`�ܕ���~GFvKk_�m>�~1kM7�[7�/X�5�<^��!�B�+���͗���鰎C�6�d�)�����e"_��4�?|�u�ZⰟ�G��n�e�s����!�3lp�C��E{��b!��T����vS�?���Νha��MJ% �W�U�U$���O��̉�l��&��r��S`������ɘ���Pʀ.�ɑMDh����a�Y�C¤�C&�q'oL���������+���#�|c��"{|���ѣ�!]�؛��,[MMo�K���~�� ���C�"H �u>�}QO������"��b�1L�D�\�*ZaVl�~K�Kq�`h��9c1) �ʏQ������=蘱�C~����B}�W5V��Z��hV�a!U��zG7�ɹXTͅ6��x�ጞ��<���K��r�;TV5�o.y�w��4�Y}��yQJՍ�{�^(�r�#�����UD�����m]���;q�-r|�=J��אU5����	o�WdT��8���O5�B/AR�4a��b�t5	3��\f���:������2y=y?N����Mb�N�t��N�����
�)C�h��y��e��p��I����	ѱ��S�ҥ���
Y '�&�T�4��3>�Z[�@����e�ǽz~@I�C��D�wMBQ�v��?HB�pސ���#� $I}�yĳ�/����d��>wa��lP���F�7�ݔ������}��i��UӤ���+X��zoذ	��[������"���h�4ˊ�-u�&n{�ɨ�Zº�PN(� *9�s`;�8�Pe�7�e�V��N/Ғq��ִ��@���oEM�����˯�C��������4<ɬ�����Q�HṸ z	���uÿH��ЇY��]��%��e�"';��yk7o�}Oطg��V�0Z�D��+a�v��e�d7(���A՝�[B8� hL\A�e� 	e`jR˹���g��T�0�w/^&a�y�VAo������R���p�"�Nc5ӥN�Ͷ]h(mp�fn�f�ҘѿQ�.E���l{��<����^]5e�n������nɑ�;w��V
�y��0`d	�d��(�Ȃ�w�l��h$���� x���3˃�I��K#d�'zI�$��|�u�ԛZy�o&en���+5��c4ݚ��4���^)�@#���K�0��$���8���f��
��L6���'�
���u��dܠ�����}��oR\�9���.��9d��`P�V�^\|q�|A��&�	/EP��T�@{�%b.�;���z�tbRQ�[��W�]&_�ŧK=�ݢ����4�}K)��a<��p�;F �i�Vm�e��]%�U�|��ӾA�b�����m��ċ��\"��$�Ȝ�X������)�E�'��4(O�1��n�%�bt���9}vd.~��2�%WFH��q��1�y�_\d�+-
��[�y�Y��!�r���k*�A�Z-X���u�]����˛��l��덲qC��J2�O������8'��[|�l���a�/8#Z�&StY��CH{Q�[�ܳ�Wʝt=�<�iCC���{��(�C��bf��뛶�~��Ӭvi�y?�es����Z�{r������ϔEm� �����a6�;�M�$���ө�ʅ��z����'��Zv�x�
�Z�E�B�J�����m��>�����ix��Z��<-�\8t	����Z�;�p��x��b;���&��B����*�ء4 [ɴ�h��Of������!�r�q�դ�#�d?zX�]���OvMk}�W���Pf��$N[y�z&���7����\Ģ
�(֮�����<`9�pb�+y�����NI��7#�m|�԰f��g�E�#��qۗ*�W ���l�9�~`��x)�f�-���#*`�Fw-��J���������*��A�F���Fٝ�i����g�5r�.�u�,%O
��a�"q�n_���B�O��xT,���,MU���*��ۜ�-��C�@@�ΰ�g>O$����F:��6/K4���*�mtWjD���pG �4����F�券�J!%��i(���x���?rU6*�H+�tJg��s@ti�����&\i��a;^4���=���ku��H�D"��K꽷Hy$?�?!$�w��
!R1/�
z��j"��э�T��R����VxQm�50���cѾL��ŗ�K_!x3�J�w1k���#�E�\�$��Q��W�݂�C����,Q��L�΀��|x�"~��V�Q ��ۼ�I�wq�m���-F(���G�������(�>܈�V�RGWA��FI#:i�9,�rM�����[�8��lR�R)(|�@��8��8j*?�#е����ד�;ZI�Z��b?�����@�U�;J��C���4#+q�ጃ��֥^N]��vYf�^⪫{ÀB�%�R�(������7���ۼgyG8�ݯ��%��L�P�"�t偅�"YHE�����\��ʑ�?�$�/�:}�*L%����3W��0��A��^�p���wO�*�?���)��`s�Ъc��뾍�9C
HOO�\'�C�=3`$�)W0�_���'nՕ�i$������d��>�l[�D�1�Ҙ���h�e��ڄ������<���a�072���8�>J(�"�l]���!9^�`���/�� ۞�]ͣܪ�&��:�/^��d�c=LV�z�k����AE�˞��8����%V.]��n�Υp�U��FA�̷R�Oƣԥf\�i.�5k\�:���|���a��I^��ȰmL
�i!�\#��}y�;��&ʅ�xm*@z4ab-jhț]^�sX��z�b���:��W?e�m�D�keb_��ޕaj6��Z>�,θ�����4
:zrA ;˿���=��(�MN���|W���Y�����]�JV�J�B<�,M��|��������}��1eպ_��Am��RSz�2�v��I&�[>��B�'5^`��>�Q�>s��r�2�G���.Q����ԩgB̊I�~V��+R�l|����o��e����oM��a�7��F��>Ӱ��}
O�ŠN����,(s󐍱[�Na&n+̳2��|��ʷ�L���"r�-�-1�0����;��f(�\�|( @�i����*� T�bFT��Cz�t������1�k�zgiZ��O���t)�&���r<:n�,��
5-�t�B\��t�p~.�@H�;��P����W�폢dyM���9�.J�_����s�B�jE[�ƪ��@I�R��_�M�J��ԭ�?_q�[z{�Ì(݄�4^]>QIܲ��]�*�u�t�5����l�1p����#��n�	4��`�1�H&?�$�^��T�&S���ZYj�m?O,9 ���y��@9
>��5�J�$a�#N�8��8�Xx$�8Q�
��Sw`�,AQ�Z2���Jc5<x��8�7�MVf
�d ޑJn�Ʉ�A>�4ފ�4r��M��?�btH��u>7 ��f��a�]���L��փD��|��TI���0����fV>)��*�ߚb��Z����L��1G�x�TZ�aiܥM0x�y``d�̦)����Q��.�Jb�o'�@,8�A:%D��)�,5X�ugj<:�nP?GN:�5ˢ�\���U�daq���D��tn�qv��HҮ�lD�O=m���5��)����������琭����[.P�KxeL�p�B�+�����a�V��V���c���y���+�6q�Fփ������۬[��7�s�m��#,�D8�J�6QP����a�K��x3��x�V��n��S��1�.{M�g��IQ�>��ハ�fÛ�Y�sL����Z�K]-zG��v���O2Z|���y尗��1�>'��k1�a�&"�A(F9�y�N���\�d	V�Rg��+oo��H�9�l�߅���(�(]kC�p{ ��1��T���c�ށ�El{F#ʀ%�&�W.I~0�gQY7����"v���	ma��Y�B����(�8QdN�u��]��;e��g�ŝ���<�\�%���{"ԅ��	+ ���L|	����SH��Ku_�� ���(9��RpBK����K�����k� �:�3����{����a��l�!��s���t|!�&t�$��.��2E����=0��:��ѷ]�L8s|~�}�0�u^���Q��Ms�6V8�6 �8�w��}RP�Cć� ��E�7<���r�V��tsy�g"��d���f4 �������W�y"/�g֥S�hv�5S�CBl- �T��kr��Wn���E���j��7����.���>�-���[���{�([Yw�m
�״bP;����;�g���ێ4��3���6<�>��0+Y��Þt렬<�2���.����D�9W��a:�ez�^$9��1@�)�C� s'�����q ʒ��|t�,�lJ�6*�Tޔr�D�.��?��8�h�����XQ����e���TJ>���+f�	�2��NTy����%��|2,iE���x	��M%��VC��o�1����/�`�#kn���#	�H�:9&��]u�(�5��ƈ�������%ݟ=��o�� �������œ��s��3��m%G�X6�0+�h������Ѿ2���i��8V�pK^�·*sO�V���	��x�/����(1!�Bo�μ��˸0	����;E:o��nh��͒��q�3�m�4ީpy9�a*i�n�<+�S>W�*<����L.�,���Q���Pdݜf�����rU�M}ds���C)=H&8�(��AN�O=؂�3�^�O��f�ΘӃ��2-V�3/���.�ۿKs�l6e��D����J�Pu�1٥�a��=@�5� q�Y����ѢW��J�"�@*Z0N�Qrf�f#�!/��m��ѳ��.����GI%pgus�񝹈�l���.L��S*	'C�+���pw�e�[��"*��\'^�62�x�jA�*�y̳�E޷u�V�,[,N��z9�͡@,��K`ܧ؃�D��.������ᩘl�ӱ�v,�j</<�XG�ٍD�ϟ��^��'�2����v�Ilf?X��&�s�䨁kg8�g�b?�_�q�x���&Oh��"���3W����/����U神k^$I�����W�	�0	�YC��0n���dq���p����������!���0{ق�<.y)�NE�6A}��P#�e� }����ڴ1��x���,#��[q<���$������xP5���L=d#��8�aE_7�q����KvS�������b�W/ެl�:_SLχsV�pC�Η���$ks�a@���WRJLo�90��k��(�s_˞á��tz52&��o�F�""�>�����ݪ�>K��| UP�`K�ܽ�s=�}%L$EJq�XaƦ��_K͎IX=��\�_���N���M��"��|�纒�z�=�e�F4����/�x�RO�Dk���NQD~���^�_- @����ur��?��T.�Kva;3�R*�A11��f��%���4�a��Ņ-��z��I�]&,~l���9,�n�J	!'�Z`>�}k/��M��t�(�R*�J6��9�2��֛�pe�B:��-�6�iW���]va�NIB��*K���?Dޑhֿ��4 �,6匈��>�Df����u�����=F�ڸ��B	c��cNc�R�\�=P�xT]zR�j2�ܱWlKDRh�w�q��g�t�q�L��&���b��5� -��D*P/o��츞i�a>uÔ|O�ꔾ�U�U�:Lc����誸�Ϊ=��l���tJ��`�T����#�~9�y�
�Kq>0�RhS�TE�4�ھ�<���m~�\ޢX��w��~�L�͉Z8#��3>K�;�Z�lώ��6�YM��5`�D5G:�ӽ�F����l��[������5�Nݟt����4�Wr�-����#��H�{l�+E������P��P��<t�8۬i3�F��
���
OԿ�6�)�T^���:���K��� �f>���_��)�����J=	{�>h�"��cT���b3	��$��;����6��p$%�����_�ȃ��u�&�:�R��62�����d���p����D��kF]U���.����U�������R��~H�{�G�m@_��0S׬\I�w �N���-��/x��߀J��=�2��� ~a���=̬��b�@�!k��es��*t_��(��H��½����G�Y�j��It'�Ö�g���Z�"#x[&$&ա��փ�ƅhXpľ�����Y2[	�y�k�"�_Km5͐���(^��>�����9�>���&�!ڪ\����z�*�be�G� �j�o+����2~>5l[��U��nSϣ���@�cyu/V�/�q��T�1�T^�oToP/k��k1��^��}:�C�r��G���p';�!}&Y�yG����R����D{�/��0#������{��Uz��RȮ�&T��]��1���?��l*��%;����׽�Kc~��ޔ� (ĢӓDŴ��m���G@|M>*?�����4�Av�)ۉ���A���c������2��\2���vǆg廿A���D[v� g���X{dpb�uhD0H,i^<�53����C��8�Re�`˘f@;��%��w�$M��x�R *V�W8�.����y0?)�>�̗8<�=�"��y��ZX���¸`�?,�qj�����X��)��=��Tϵȓj��[0�֐"�ǶN`�ܩz��w�M�c]3�$d�h������܋:�������5�SN}���3���g7,;���;C���(��@Ҍ�Ǣ��$���5���,�����DR�	8�rڳ���J.TT����t5������c�ׯݒP�-���� ��~x��O
�α�x(����J��-E��c��iϯ�|�,�et�I��X��U2�wi�i/�v)$���s��c=6��֭ޜ敃����=�M�޺BN�3��qCe�䳡������f+qRi��fi���g��p=�S{��>o����Ga�22wr�M�"�r!$�cۖ^����EkC<�l�(�O���!�X��x`����j�������'U&E��Kx0��&�c��a��<�bÂ�-�XB����e��q Q�O��{��m��R�������%�Z�����K,�~_�fH��ψ��h� y�����r�C,݈E�WfT9U��ew�����J���������Z�չFBĜFd�WJ�<z�=�em����<t������8j�ה
lڶ~'�ϗ[eR���;�@��sP���^_�!�7�������s�D����
�ʟ/�<�E��eAd��y�3Q��C���2����yX�z��# Ĕmb)q�k��6f$]}��1�Q��W��u��Y�-�N��@�>��������S�-Z��cyJ��J￈�W���&t[�2$q�mS��J	�/	�q�Siɡx�9�b�zV�7���� �m�` ��4�d��_Z���|o������R����cE������w����$�w����w�x}��]��l�7���]����t������䡂2�^o�bR�9x������8����ul�N��4!xo�+�|{J�=�2�{ŭ�lMٕ�/3�z$�菗N4"+Û����N�3��҂��}����(Ev���8?�S�3W�k_�(и��%�� ��y�o�)
�I������9|��_���Ǆ+����x	���RZj�4+�{�kl���g9�1I1�w�����QF�1�Y�
J�1����D%����QG0��	�&p� i�������f���-�,=�
pi�W��E1��yr�K��`��C����#����K�Q���������ޮ9���Q�xsu����yv�'��Zd�W���Z����g����?�ګ��X3�7c�C+Hu#kA��"���LO�ܴ<kM��@�o�������ÝO�FI�J\�M�a
j[�o�A�V��L1���4fn'�b�����M�o�-�������p:�(�����z.o4z�d2�N��V|/6��kO�P�LZ��;rM��3��|�K�j��n��eFB���?�5�~9*];gЉ�x�� ��	`�%CH'`B�c{�����0�Z�FUH��~�[�#���<�,����7L�h��-�������S ��:��ÅuE {{�׉�<�^<u�6}�[k�ma��.�m����HzY�A�Ԩk<��7�ƞj%�w�?3ÿ�KֹR:l���_�_��*����э���*�x��	(�dfN�GKx0�p��g �|b����/�j2�M>���Ĉ��6GK5��f�U6���V��=�r��z�<܍�6<"A�Q����a�?�y������_DJV�x��&E#
9�>�����U�ݦu�Y�7��=�7��-�/�O	f�f���\�� ����W�Q�
��#�/mD.]��2U_nq�)���~7�\���\�ȣ����K���b�MưZ�(�&P49�ɮ��X�>��6����ޘ���"����!4v(Ƒ&Vd�Lh""j�5�p_��9Έ�/���	B�AHS���:�9jw�yN��̲�*oP�e{�$1��x��c�ϻ�_����W�Xt=`����T��h(�|Z�F��xo�^�"�V9Puf�w�U��׼����b��p.c�c��h�_�D3f4���� �X9���hdz��%(�����Qk�ř�A�S���f�Sa]%��_�L#B��y���47��6���蜪�ʹ����S�;B�(�/8���f3c�4�2Q&NsZ��t�։H�ݵ�.QA����(����$�xC9���.��؟V���%�o����U?]���+�q��$KaQR�E����GTf��s�@E�;��Kω1�K��-E�f*>Do����\[V_Øl3jI�D��{|�,"���+R��=j7l�� ���>��~�FS6���$��7x��8�34��ס�l'bU��m&ٜvFa\�ޅj�8{+���A�(����a�{'�Өء�Bt�Bs���J��JY��*U�M�7}�3�싙���0�xF=ô٦���e���bHH��ص�M梷s��90)N2�Ev�������=s�Be
���*-f3��k�@.�{a;����rq�U_9V������{��&�d�������(�obr�ds?�|ĖK�A4�X���G�oi�I	���}��� ݌��Ûa�n���N�����QU惩#�� ���-s�!7�Q4AhEl�<�N���u_���<��8�h�/8�E���5��l<�S��ӍY"3��ԘD���t�
�������=	t� *��� ,��H�ڢW�7ي�������
Ho9)&���:*��B�%q��1�:��Ĳ�Bo=�!�c����0IA�~	C�,�S��cD���c��_��$p�C�鞶��m�Ͻ7�>c���[}���P/xDޢ�)�j��%	ݵ_j�����O
ܽ�ա��FD�Ǖ0 w�e��D��
O�&B5�s�%.:f�5� �ؤ���9���]�<������>��H(���O*��e�{�� H�u���eNxC&�t$���k�*�uY��	`t(��	}�B�(cp1���7oE+j�Xx�7c�\r��`:��O�<+���5f��C�t`������V�=3��X�)E��;���2����a�>�r1����,�Զ�����#4�
�Y�f�BY��Ç[�WX�4@g����b��=|����LbO0�'�K'��G�³s΋>�N�����Z*���瀠Un�|������(�2M�!��B��t��*}����䩴CDLF���{!<���͊�4�5�W6;��ǖ@-T7�Sӎ�m� ��QW����j#R��$2Zô�n(�ɑ/�D���Y��)U�fV!�w�C~��B{9��@r��));WtsMZx|�L���+
�k���b�Z�$�ۅ���w��Gb����u?��ȶ�����* ^f�J�!�v�m��s��$�;ֺ�8~���%[="	,>0N�J~���_F"ց�35"��%?�R*����,�[Ԇ=���E�K`M�0�w/G��4š<0�Wk����]sڍ�����ծ>���<�����<��G��b���f��m3�PN�&GuȐ�������ׂ�>�7�*RP{��	8��2�ͯuǕ�ϫ��BcV}�2��0����Q�r��¸�ϗ������l/5��CΧ}E��e�M��v��@���r������)�@��(�Dh�B����P+gQ��	����Wk�&��)MCx�����\<���:nh��U�m�:r�X_�!R2IFld���m��v�iv~M��Q�k�a�@՛��5�7:�B��|BǌP���R��H �GdZ�rP�8b��j�IZm9�!A2_�({S�,΂�a�[�` k{jd�R�-��z��c��K�-����ߠ���lݣ̕vDĘ��E�k��C]�_d�� �%z$�'�Mً�Rk�E��`/��]�r�.~��
_�3�>�A�������mv�_��G�L|�T��ũ��(���H�b��\���FJ���]=�-��ʈ/�f361D"����(��}*�L��q�y�/#{o��-U>aR���$G�Gi�7��h�v�ۍ�g`���I�/��(�3ij����4�Y���v����#}��'ӕә]d����ƣ�c�������}��U��R���ye�.�*c�vQ=�>��x '.�<�w"U���(�����-j��
*���(si�g7~�Gj�ɨ����
�����(��䦓���7Zٖw
�I����XD�T��!�b^��W���I���UeH�}�?pC�<��,v&��0������A�aP"]h����$���C!���`�gIɖG��v(�>����`�t�2t%��h��`����p�7�?���I�;���2�UrB�Y�|��S����]���̪4�ûQ��(�d�i[�?pNy��`3��p��K�1�d7�]�I�/����+M�������h�o�[�f�Nr�5

���<�7d_b��_�%������&��"=#^�'}#��}�z�뇓It�R����驪��r��1��g�G�G~�����N�or�W���!���-Z�)L��\9�:Al����2�6��Y��y�<W'��c;�����=�W��E��J腧r���^��u��[�brI����XP��7�!��=E�9�2F��L�6[<���z�B����+��%��j��養	�^��q�� ��f��~��"��{|�_�v������dto�KПɆ��`��U�rsWˏqQ�3�PZ���+e�����	T� �\S9X�%����OZ�v-��2��f��s���A ���@ፖ\g������b+���;RF��(������.��Zz�p6��� ׼�V��W��C�*���	R��W�E����n�a�x�;\����f�'˗�b����b�gd����{A��P(V��m1�g��nP�Y�a'T�?�K~߽�si9�F��BN�9umE	�������EP�B%��@R����o~��%!h�T����>�w����䶭��t�@S�,�a3��i�}�iW�<s� ����֚�K��>����<8�ھ��Z�V,�Ȥ��L7K~3���-@�	��yX���$*]m�헽s�!��W�^���yDIN�u*RL����t�'�)��TiE#�^��@�L�Pe�[a�x	,ެ~����u����C��R&���\X�憣�/Q�`�泷J�X~� �..Y@'"�UnF�>�8�M�\�%�z1���	�G�MT��>+C�#ڇf�6qo�b��bO��	��g�A�y�n Q���t��u��Ȍ6 U�}Z��!Fm��z���҇�-x���-?+#8vFr��w�f��mU�e���M_ژbu�]��3�"ӚK��?`qT{껳�H�$�-��C�����4-����p��nY��)U�3���� ����Y$�d��.�7��(��,)�P�c�4%g��İ�s���Y���mrP��6rp����XS{0�ؖb1�&�{ -=X_?���W�<���5�J��!��b`"P�;�x���=��� ��3�&\��< ��̚��0�LW��|O��f\�M���b9jM!�w����ɴ�$A����v��eՙ�sZ�1�4�oQrHĜߗC��s(�Q�E����\I�@G��0�� �"�㨌4�4C1��ۉ�" �vm�#�p�'�ᷧ��glxYu����!e������̽�5ޠ����� �O�GKd��Kvw�P~-,��i u~$��k^O+���(KY�I�;���c^��ׁ�����`���7��x��"�=̑�j�\g� O�!Ko_V�N�\�!��S� 'xa}�@�Q�Hߺ�9�� ��8���y��%&��o9�3!�M��To�ka�7 �D�>�)�k*�>�N�v��e�g��AD��5f��޽DJ����(5t�m�5�y*��n`ݭ%�$:�qGP�|�ݫ�������Q3�ʧ�o���e��(7����8�HEXt$ٞ�6C-�ĕ�S��=GM��ʡ_��h�>�'���k���+n^��:�5j�
6ى#�E����k	A�	�K��� �:���4�yPǃ#�+ܦ�?A�;�����3|�kj�s�� �g�D�Rx�2�����iἭc���t�X��PDAX%�ę������ݸ�ٲR+�׮g:��P��{�L�v
��U5��1�=|r&�L���R���EO��4|e�[�LA�'}�+h�%Iq���?���Md��(:�����`O�l�v���,����*����'f6��PW֐}��E=���MN{��V�"�y��Xb�tA��z����)�@��r=�D|f#��eA
���̟�����-7oe����3���YT��\�6�5�n���Y�ˬ�o����i�����]>�$r���B�l�ӫqxn�+�}�F�΅KV��B�8=52�d�=��7�Ϫ1�<Ҕ�������~�^tdq'Mpf���ԪX^��H��䍅�q�r�d�ۀ�_�̼�5I��x\>K��曶��P�(u�m�mg1���,M
�3a�] ުT��V-��',���Ei�E�fH�!��%����Fb��]qjf!�i���/��	c�o����|��K�[�>�L��i�&F��>�I���;��������}�b�����O��Rt"�BJ�#�3�C']��� m����B��v� oY4��#�b��R'��/�ʣ#�D��* �d�����3-���¤�H��T`j�V`�o���r�J�v=�3����1/�O�e��-��?�ܠ"�T��o�C�[c�P��֭KP�;)=�a,�!
�~9ǳ�j����ۓ1U6��*�h�����Vު�ife��x�GjSC[��il�镸8�?*����@��\j�y,���!�֒I7�| �2/�����7�r�Q�_G�TJW3�՞�=��R����i�݂�;
�l<O���7����"v���*�o/`�6B2AD����A؄�n}� �n-u[��v���O������Ot#`���dڵ��tm��x�Vo�)@2M���|D(�j�y�A����)Xh'���|�ﳌ����(@�j�gW�1��ʵ��|�AH@�ո�5}��F�F�='�{�����t�Bk�P�[}zN��s���wx��ݱQ�Q1&���!�07�u�,8Q���y;a�n����g�����K�G�ar4q	��8+��`�v��U�No!����`�'�sw�,��]~�y��W�b=�I�2��G��F��➱F����I��s}��"?V�E��ゐ�$���33(`��y#�Oq-��bȯ��R8�͕�H}W�bu74{5x�_ڬ�.�[� �l�!�O{{x`�z�UO���LT(9�|P��Ο��z�D;����c�j�ZF��3��;��F��r-T;�BQK��W!��zX��^ֳ���Ƌ!�*��>�O�"�a6��g!a�Ua���Ej��N��stwNY�7�X�ҋ���G�������J�e",/z���J�EQ��3x��/:�:^��@�6����O��7��� ��k���8d���4xt)x�;�`� ��[�9�?���4Zk]G�-M��qR7��*)���	z����pz����KA��R�<�V�C��pC⛆�K�%�;����<(8F��R�L�!�Djb;g�a�ʳ�;reb�(�A�y���^�x=f�"ۆ�4d1c^vR��C|BU�w��A�tl|>�� Ո	�e�#)��\;�H͍P
�`Uo]/,췵��}Ν1l1��Kg�3]G{ �C����Z�hYa��7�T0���֍��S�Y�U�V�(�IZ�&|<J�q���n ���ͪ�����9q�A�X���ґ�m�z���pA#�uw�T)市�H+p�K�x����h�oњX��C�H7 |�g�f׭���ţ�I����ڏ���8r07R��)��]ϋ�x[P�#�p_T��.~Xj�!�{G��-��J,S(�UT�a��Uc��$��<Y��V�د�?�����Y��-r��'i�US���V}�!WYpI�2�SB~��b��w����[�dg�ٖH%�����R��8]V��T�<���̔5�P��eMũpF9��#h0��>j�9���ڽaͼ����e��R�ݾ;����P��3༦"�d���+ɚ	֏v���ZT��Z�j�x��d��ۦ��l�l��,���Ĵ!&yM�;��4O�1���1g��/�E#�1M���$ ���bo��H<Kx�v�~����l��f��vK��f�k��鞒���8w�s��(�^ʹ~��������
J�L	yJ��=i�%HUH�#?�[�K7�-�
�L@#�A=!Kj�9�Db�-N����B�d ��{��9��`M�B�7�L$"+�_\ؑ��/G�9%�^�-�,�}�P����K�j�/�"e�����I�H�%8.Nv�41�U���m�>���B���d<b�����Z-&fU�6��7ID�{F��?X7�%���~��8��=*V�N��~cc�ԛsl����֨��۬�#q8~�^��lZ4��ҳ�\����<��l���e�Dv�%%&!Auh+����J�M�ɿ�8�ؤT/�Ǉ�Vj�4��,�r�U=��(�X������w�����a�6��ŀ�	�\��,�mI�DJ�$H�h�L�}%!�#�E��뙆D���E�Q��I�1�X���VX�:�?��f��x��2���X�dhd��A���G���Tnx|����`b���v�2c�0�#s���6�S�����NOsݴ�e��h�a�����ğ��NU_Oć���Kf��s=���7�mN���%� F���3��>˒B�b�J����S?������J�h����\XR0�m�������u'�T���9���KŪ���!t�e%4A��2R�ƉGCwhG�|�l��Ş=W�/��,)������?�kPI'!D6u�)0ZK,�[���{j%6�I0��W���@�T[~?�<OL��P�l{P+T�s�D�jP��H#"-]��^R	C�"[掄�c-����u+��xp
']ߧ��p�	��h9�+��g:c0�5A�8'M�YA�L;�����X]I��˔C�oq"rZ�Ec.��\��{���aD6;��m��@�;X������<<�ΣШ_�����u)1f{Q{��0������֖��O��d���LQ����[ ������A��*l�M;r��.�5�;���*�Dz��<_�C����ʣ�e���Y��յ��F�5_ŖK)b[0�[é�e*i�������3��D<��DWho��F��T�Ĩh���!ݰ�M�[4��Y��|9��+�]$�~����Ii�T	��`�M��Ȑ�<���TN�l�s���귘Z��_C�}����1�C���H� ��y e[�K�Y-EfѬ�%��m����uͧ�e瓝˛И[��1��Q�0�fu�I#0����}X�	8�+y��=Xg��ڥ<�8�pR��E�0���X8V�(��~�O�u����@�ߐl&�G��s�)�yqS�z�?�qSQG��_�"8���61p��3	y�?Fm�B8��Hn2څ�Rg��h��h%�K`�Y'��V�iX׫�H���c�l��Ǉ�l2��ƳT�죐�eCL+�!��I؍ܼ��Xj&��Y��&�n�ՙ�	�]H ~��_���]�KD�vq_��&�ǩYM; "��v�`�B�e�AD�Z�ݎ&�mQ�g��_�r D��S�X�u�Zy��V�C���'�q���?.	��1��8Έԕ��JD��S�O*K�wר����2WS[����4LY.����2_� �*��G�bnκ�+�w�G�^�m@恩z�H������&���G\+dR\`F�NT��S�����qh|4y0�Z�o�R��;�3�6%�Fuq�o���`M_9�<���#x�Z+��oa���u��l�]��{}L�'Z @q�­m���(佫5=�f\9�q�@%@����bƝC�Gǂ�ic��B�F%e�R�ɾ�{.�-w�Ǎ `�w����6Y�_�0�<Z<���ڂ�hj&/B@���؏�L>� �[���5�O�hoc����y�P�*:?1�9èR)�Cc�i?w_T:S�ɹ��f�! m�xN�ҁ]�CG��'��*��TPё:�Eټ���`���E�{W赡���P�e�4����~Ib(ɘ���}2���k�������؈��X�v;�R�4��u�f>]��x���5)�l����ra��2���v�����_���M9w@1�s��
�9m�E����	 _ǽޮ>p=�Q��az1��\��R��%>}�� �4ۦ"�������<Y��GU���m
��P��$��Fza5ʗs9lEG�G@�|�T���`��hیF��6is�z�x��3�������t����3<�m� �)�E�Ƒ�^}�؂4�7/�����'�Z���v��	���fcqSתk�%5^
�Æd�kz�OL�w�$e�uG2�<.���(�j�QΝK�����^�S������\Z�t�Ż2�W;?��b���9j�{i9'ǒH��=�h�t�C�Ƹ�F9N�O�a�s�g1�u��5�(�k������9v .�I?�������g8Jf5!�y^��ok�+�Yw#�����J=̵ե;o�I�ϯH�ߟ�qL���6������F�G$31c���}��y��q�g�n�@ 1�ɝ��+z L^�X);F����,ĻD�lq��0>vֆ��<jŭI���-�@��Z���d�E��:j����iD��S��o��JKj(�w��["�E5�����l
�I5��%���*PJ���Q�S�����>� ���4�dh�)Q1�=:�[������ �;^��"y��I05��iD�.N
�-ǒl�g�������P��do �_{70�cm4$�޻�ayK�	3��-�5��5b�_��B�k���[ǵ�~�
|��%ӊjR����C'�x򝲊��7p����Vh'��U��nhr/�Ag=�������r0�H����1��0�� >P���g3ힷ �P�|��Vl��JY��,e+�o�J}a���5�إW����?ra����V[CN�j���U+�^��C�j���~C1��Z�4\�>�Ė�XZ�s�$m.�Eޅ�E��.��)��G6��׈����v�YnL�����T�HR��?9<�nd�t����tS�V~�0�A>���V��L�j�� 3*t�&��}�eɿ�fa�S��
��cE�4N�bZ" �O��SBCR�8�c�m��/+�/����H� \��n��[�WTv�3&��w>�LZT3��X�=�Z�RQ[�xc�>V{ۅ��NG_me�[[�������NM��^��6ᢌ�j�se닥�n�@��|�e�?����Od�)��ΕY�6�$�	�C�X�r�P)�~TS)Q�]@u�;��+��A�$~^is��Ã}�
�F&��4!T-؈g%����p��r���f���2��"�np(�,���k�xk'B7��������UJ���Z�"&�~bZ�N��H�h)��S����+�2��I=�?e>�\p�����4�(�/)����(���#{F�b����)�3�'\��oM뜃�i�؝�B��$��ME��+dh��yIT���fӂ������}����r�lZ��jMi	��(���-Y8-���� -�cVz �i��f�R��ì�*�3�_��	l�8>��pt��,�DP���Փ+Lo���)7}5�*���Hb#����T�)W��� T�IC�~r��ͻ��,>�ڲy��Z�ٸd<æ���d��Qr�3�슚�C~o�x+����k�^{���Ъ��c�F����ߩT����~]*�@0pDc���r+������.:Y�z��,8����B f���r�ΫQ<�T�"}tv���(��^�b;)b�tPS�ɸ���b�NN���ු�~U:_p��k����C�ԨMl�N]u#��=��»��!y���T)aPƏl��TxŸd�'�Q���z��f�t*�X��}Ҋ�e�0o��%��L�*Jd=�Ŏʕ���^���,�b��%v�݁�]-��T������iǟ�n,�"k�1�M�P:�Kg22.qp��i��r��� 
��Bq,ΆYE����}R
�!�����4i�	�_%+��<a쐩�y�e7�F�[R��H�R(��2 �8k#���W�G\!�v��z�|xN���o~���t�p�m�$T
��Ŭ�M�-u�Mj�u%���&�7�_;�E�.H.�1�7�\+�%����l&��6�"ޚ2�wZ>@��t��v���GaNNy)� �9�؎p#�⇕u�3�/���{�� @�%��H;<rMD΃���ChQ�(�5�D��@v7�T4xB!��oC�#PX�6̭:H���T����f��N��q���)<Z.�x�p1�%�_|���������mk���{"{?u�,f5{�����M�sV
;S����4��f<���lv�w�g�{�Hh	ۂ[NAp�wA��#��r:u�Fa� P�z.�H�1�8�aq��v�9f^�����A��z✟$�����5L�x���w<��qxN��'׿>���ʢ؇��A}QM>����@��s)�Ճk������/��ao:����<H��W����D��Is:��x,}�PB���S$��)�v��皱N_"l�*�D��4N"|XP�S�w������}��/��
|�6�~M3���f�����Ҫ���ɵ������䋂Ǻpf�y�g�]cx��!cr5\pwFPI���sq72��7(��WpQP�Ľ�㕉����3���T��~_Db��(��PheL3_3ӳ-�Hg*lPa	�;m�R6ɳ���YR!�5���7<�'�����c�hֻ.��4&.��>v'�����g�_V�K�@�R��>�c���\AF���Es�P�J��sM��qf{㵚Gg!۟Ŗ�.,���5>^z���_��J���i���⚍���b�L���U����A����pH��z�W�U~����iQ���ϵ�x碪f�>��=����R�2��_���M�&>����� BL$��+��i!�����4���f*�}d�����E-���|S[�����}F7�<P���s�9���88�U��vE��i���Î<�M��yn݉v��Y'��7y���)W�4�_�
N�#���1a)��ՎCA5`�	�]i�V�� �4h�[L��S�[�t�����ݷ���Gc�?��^��Pq�OF/+�8��q���,��O,T�6x�����C��t7�}��PZ������*���Y��)�Zi��6�nz�6T@�G��0�!�= (�q�T)c�q�p�'�-z�/$z��J΂Z��Ё����
��އ��W8�!&T�M�Qyb/ɷ��-�^�g(�u#�7�>p��g8�CA�̚Q�pw٤���bN��[�ME׬0�5f'S\GH��Ѡ��R%�J�0���[D����v�R|�ᰜ�.�w�cf�ʮ'�!�4n	@���hO�1�l��n��ԡ҅J�Z,�£�=��K�0��g�N6I i�Ebm�{�;Q��{#!n��>g�l�t������rd߂����m�`*V��!�š�c�2"���K�]ho^�t�ow��GJ@�~�rw.��l� ˦�QaD���� �4�π�Y�
� ��8�(�%َ,����/�UuX7oc�/�М�4���/�H]��M��Q�3�d#-����F�������j̥n3q��%E��m�[�L���ޏos�U��z�(��a��I;]�3aYb^#�D��R�ᐢ@* ��"�Q�*V��N��Ȅ[1|IZC�0�8����0¼ ﵐۖ�j�ފdsF�_peh{o��G��e|�I�}]V�5EöZ��@��SO4��� Y����������H<53r
S���v�����������g=�.��u��������Y& ��@�O���C��>�:��9�T�(Kcօ--�w����
tj�Xs���*���~�;x�z��)�!����*{���2�-����xc5w��r�D�B�S�h�(:�!i	�x�w��+�sgZ1.5� H¢o�o:��B����`Ǟ.�$,}���I��>���7`k�j�7��ae�hk?�� k��2t�h#�Uf�3� 5��m��v�Ҳ�F'鉫�T��T"�H?q|���O7���g/�qzi5��,�.u0��&C*s�E�C��ad!:ѻoQ���������7���2:�B�����- ���l����VO������I8y
�����Q����o8B�����r�'9��S�0��}�F4��D��.����./ʃ��������_�J��i����^�[�=RNx&���k���t	Q]_niB��tԑI=�LǊ�TFO�dD,��	�J�y������".{7�];D!i���#�K����ֵi�1�?�W�eW�I�U/�|t�6���-��9�F	��#�������*��i�ڈI��;��M��U��������QpMs��W N�bQr�?*�+��dL97<��P�/Ts��4-2a�˥;S+C��dd�I��ДP��jMe�S�:�h�������[L�ԙ��ҳ�M���=�|`]�y�i�����Q�6�?��,�k_��c��?ǘ�.�����9{dЈ�FMG�lg����#��O��1c�C��]X����կl%$�/���5��^4�׻�\���� ��X'�v�6�̖}��}�
������`�h?�.k���ra��77�\����FYI�������gsl��]}*7{���}�RB]���)���t��s-c�� 2�t�m�E9Av�]v���RC+�Z����B�1Úh`�%�M3H'F�<|?�Y��`ۍ:j��yaGr��W1��bO[<'�B21(]�Lf`j���ͻ7}�����B�^o��9%"�ذR��m�̜���8L���W�n����Y�o�nd�#�z\	�#y�8Gx"��q�7�HO���_ͨ��r�����Sr�(�ݾ�
�X�]A�}�1H��-ො1<+ܾ�ysQ�l*r!��R|�F>kff��8��9dY�mP�"�6gP��z�f��dϖ��]N���3ډ�ɐ��1�Oa�ܔ����b�kk�|k���(�1�Ԫ����<��*ʦ:���DS�:�W����(?����������1�����V'0p� �z�N"�w_�y��!��T���}�\ș�	�p��[^r���m�+B�QS���?�.��g�%��C�Eӧ�\T!�A�ݘ�=������YR�DԊ���,��]d�E*������9�L��+J%u<μc̈́��E�K4N��G;�W^��6��Z ���G)@9!�&�C���ҕ�s�N����/o�]2g�ZV��hȈC���/b�,����"sˌ�eK/P�=~�F��)�wpa�q�YDḉ��Q�^ �l��j!��cv`���Fr���'��2��OY�����&v�y����n ��t��!h/�Z0r�Ӣ�=yUU���s)�ٲ��>��\O��q�wq�/�nw�,~�ra$sVf�T4an��[���G�ʻq�����F$]bw�T�bM�J5� �e ��a�e��=�v�5g�Z}��1;� g.�댼�3F3BX�D��R�&����#�1f�N^�_���d���Ǭ�D��Љѡ�����攻�2��){�����mFr�lZ�����D�;4�_�K��+_����g:���i�(�>3�=���W4(��?'T}{7-�t8�N�OSŚ��8�e��0��bC�&$�G���z�*���u_���_d�T8��ZD'N`k4�&������^��H���T􎺁���zzYf�?�j����_,9?U�r�j�h��2���A����֮!ہ�T,�kWQA~��P�,�K.�pJ}0+X^�����C��8Ր�ۥݦ�-����8�[�wf��D>�ߜ̩��J<&������Ena����gf�nW̤���P�ub]B�CR�7��*�M��"��P}3��O�D������-}J�ԣ�S7�~0K7�F����]�ݒ��OF=ɍ����lQ���=��j�.%�6y��54����#�0<Y�^�`�"�-8]Bs�j~�#�.D���̠�8DNz�a���k h�GT��@��X�ĉ`gת�Ҷ�zpX+��"
|��ﾫ1��(�&�g �w�^�?�,A�	�*Z0��Hjh��P�����J[��,I���g��P�\��[���"O&�w.gt9J�JH����\ҝ~H�8���n@l�rC����&u���BM|�+�����܉�P6J�Sw�����'�Bm��@����$�Y���.q�˧s�P�70�)>�iL::�X�NΒ<bz����P�{��I������/ �G e�_�.0c!��(�
�_l�/���]i7��5FS��	�j<��w��C��ai��e���rZ�MFJ��JP��R����8��wR�",^:T��Wv� �w&�/([TV]X]KFc�B�y��L��N�D�*V����H(�C��������xA�Ό���M�'5�I���Mau�D�Z΀�v�";cg���u/K�RVCu�ЌOh�B�:���r������z�a��C��m"�֍��tx�1����*�><hi�]�Gh���[<�c��v�:��*���w
��]�*z�5x�eK��Po�ҭG>�!�?��%Q��{}jK�[��3K:J7�x�sd�!Ϭ� �����m���~R�Vç�cL��qv�7�.kX�)��_WH�
?\/�=�״q�0.!E�������-.�d���1R�h"�o�:\4�uL�ї����i�|ð�p̿`�v����cDQ�-���Զ����9�O͝�U{��LU��*z�W����/
���];�ę�Edc�@��c7n���!���W��� ���y�b�Z�W3C�p���Z�+dզ%t%���G��I̍����v+�,�z� �׵�5�66����(Σ�|f~R���=�׬r��*hwN�屶&���;��X�/c�+��4�[]�m�IZf��No
�6eI�$-��/��"ҁR��j��{��<X�ab��S6,��z���,:�!�N�˕�,�鮳��E����5w�Q	n��O�C�]]��*�~]m�\�� ��H�i�+�<Ο�����ʄ^�T����/x&u��S<iM/	���F�BG��]�xk����-hh��O��[Nýؠ���HW������tL�(ƾ�$�z�# �j���]�� &�>�X>�)|
�]Vz?B]@��MD��Ss�l��q�@�9�'>��'���-�������'}>���ƼA�j��U�8�����6��Q�����r���ʃjh����c���l����s�&�&�~��4�3xs����+��4��O��QbV( suj�'��?�����a��b�Fx�˷%��#~����=u!�����1�� �/� ��4�vK���{�T��Y�ٖY�HɨL*݈8��5vC��심�˝"g2�Ӓ�Z�۪-����/�r��m;�=����ɣ�=��K+}�c�2!�fw���J�P
�J��F���E�&.ϺH�"�J
���h�V,�@w�&�e�+:�߫�t��Z����Z�~6�A���!	]z{nKz���$H@�$K�t��)p�[6��t�w���!PK���Z���;e��%�jR����`n(�п��H�p��ۮtk8�����aPA$�'�6�� �w�
~_�)�;�T���#�8p�50Pq�E�籑��w��g�0���g��3\x`$&γ�f/�.��y�������r��{�u&v��P(�Da�U�0�D�~;�hMC��BA2�l4~�cA�P��+�l����"R� ]aJ�5�f]Ui�~=5�9Oi^C�(�q<�<�%�}Ug�;�$��1�*�m��Ȝ=ݝ��k�S��̮���X��w�;����Ӑr����?�O�}rp�	��M�C��J"�e�"���׽P�%�1��>VI0�la���ɠ�VF:��~���M��<�)A�ʁ��� ~|չl:\O��m��P�'/�Վ$������ ��$�5=�	���@e7��'�/<R:�Fi=��wx��Z�.��4�.����I౲ZЊjRC�@
�K&��dV�Y<T	:�������w5^�?1������Ӏ�> I��f)�����}��������z�_#�7"-��?�g�����$uf�C�*��P�7�]S\܁<в(��]�Ǵ�h�ZF�J�����"�Uu�,�P�<��i��+������́�[�Ip?�L�
7@��i�[�t�jn1fL&�C ����Ʀ�tdN��w��n���i��
L��͸���.��X��|�4%��BUmN*%���o���8��(.?�O �^�:�ڼ�}$�*S5�a�%�'�Ռ�e� |��>��5��5<5�zX�Y�x5�*4��<��#*s'ЀgⰙ�NfL*�<%j,ΰO��@%���8��!<���-��R�Q��&f��T��u�ޫ�%"�#�d��G��&��=:�Z��<��Ɍ�q\_���ƺ�A�u����z7�f�pv�b婖g�LB�ZA7�\/�:F�x1���C�C籀X��!�G��:߁V�h��K�,����۷cv�"b�=�5Ϛ/�Ho�ؒ�xrw�.P��<�+I�Q"uf+P.�s�F�řuMÂTYr�Kf)��>F��j� �e?��q���F8�9-r�"���� /��s�?�U���\�?���ԟP�B�G���\L� i(��2��%��U�.x�d�Z��~���h?'9���7���.���9��������\+�kKv�����m��/@Z@(�0�kno"��᮷���r�sB��l�_i����We]�G�[�d��v]��q`���/T�e��߫�MA��s�q��4v�Ş-�B��z,�${aFݷZ�쟎
0"滛p9�H��	��V ���>
g~(����tB�(�It�$�!�w o����mS�VL������M\�e�����\@ι� h�<1��c�`��3�e^��.�.��[�Y�)�N��'���t߈��_e�+p:Q0��3� �H���d��Jv�5-/{YQ+K����i�Զ-t~�v�kG5X��}���	��ow�h<��zX �k_^�_߿����,�ge�Yi����,0ܨk�E���SL�=a/����25�󨅇y�`qc��Ҽ��
��<PF�z�G٪nk�O���_�ScԹ�l{�NB���*��~h4ZD�N:��e:D�"�W_k-#��P���2�єl�R���<̔7,��>{}�BSX�eA�6lM�u�؟�W�&Ǳ�|�M�˰�/�ɶܗU�"�a���,�D��W���ܵ�C74��QaV�����&!�P��B�I��JX�W)`3�a�r�.��^�y����r5���(���I0f�^:./BBc��U��N�����"�ܨ�Hj��_���8�"����'�J-X��0F��%u���5��-Q����~W�D��OA�XHO�@,?_K>K�N.>G�\�$���A�Ÿ)'��h�3�")|����4���0�	@��_��I+�)���Whbm��Rm3�sqP�p��o��A��~�}���һOۂl^��|�R4��O��~�H%����El���V�b�[""W)���)}m2iM���q�x9��Ȉ��OP5�"�w'�@o��?�c(��A��8k�,���Q��"h���}` �n��{��.��=�S^��5.��5�Dn�^ ��h�$aM��!+&�F׸�=�-SD��.��n�x3��9���,0V�+��HN�z��[�1��;�u��_���<���������:���O!�EG�e�ҩ���-��~�� ;�����6�^̗�+����t��c:�bIn���[5z��x��[�:�0˓�r�k#�6|Vϟ����<��l��
bcV��m�蛛�5;e&�0`��E�ӄYhϨ�U8�G�MD�Y�98��S���"3M��ѩ�b6.Y��&~[o��[3�����ϙ�k@��V��k%��k0�L�J%�5�k�|�����7y�5@�`\6΂��3 X��]X�}x���r�J��d����AU_&D���۵�XL?�m��>&<j��K6�?|:�X��$� �~��,�~܆ʮ��"�~�D�����c!S�����TQPM�t"�3Hl�`�h�A�_���}��5�o1�?��RW:)�/��{���˧'�B�Dc]�9h����7o3���FX������Rش[��|��A���!�?�f�pt!�S��h��1�7Ix��?Tأ�*��v���uEV<�n�QO؈c�섻p��lO1����I�~qѦXd�J�޾��<�BɎ̔6Ĺ���{�2��N�M P�S�3$lhi1p�����:*3$m��"t��cJ�<\�3`��c��i� $�2�{��x>�$i�\���Q�U��*i)�cQ����h_�Z\���$�����q�;�|[��1�o�4kMJ-�f�_���˭A�}ל�&�W9}�Ͳ�h?�-�cv$�(Du�?M�̐��U��ضbC��
�ez�!�o,"p:�����P]�%�uQQ�D��8���F5e�:�f��A�PcSpLIs���z��5l�0j���j��4[$���˼X�٣|n��s�:Y�U[�⳿��6#�Ik5W�c=LƦD�"c�y%��q�޽���������l�S��5�U���)�E:������%n�;JKt�͸:���m��˚�|�����?[�`Oɾ�I����8�X�C�(�ï~����<���񌏟Jf����>�	X�[���MŮ�J���8ϿO�xa6�vʤ��W(0~�w��N3���p9i3��D��B3�<���_�e�mS�kq)Yd^���}2X�!-0n`�&jЙ-������{�r�7�����2S#�ɶ�r�bep'�3|�.Syd���\�/[�&t<u==��ZOnP3Ǿ��8�]+A��9�j$f��'�ކ�n}ܙ`�]B^	�.�Uwϓ����D}y�M�5��Y�V0�@f���%}FN��i�c綠��2���.t7���[#�(9dǖܿ�Um�o��B�ʿ���������;>`�͡-D 9�i��%k(��n8̲bO�!��`U����a���GKe�S��������q{3t0�/��` <p	�r�o�ւ>��(������典,E/Zc9�c� [|s�o#�v��Y������k��]z�I�j�V�����3@��<"_���.o2X���[x����VD�6�Z��� 6�e0l��������Q��)c��ce���#���xG�F,��u��Rn��ߩ��2�Mّ =W�����Ky��׆�8
�W��Pk�(�{ܩ�ByP\���.�iÐ"w�
�X��a���15��ǁ���[Q3M���sT7����S�`H;��)�f�4���z(�-"���)�u[�n�[�<���Z��c]<�M��S�d�E��p��nM��5�*�7d3� �K�V����JX��O"����'`���wr����썂��Aq�IAX����ţ:/I��V9ɫ� K�o�'x���r9��UD�	���W�.��[1�&WD���=>q�Ηo��E�0�pI��z�ĵ��>�,+�/�M;�Gy�\P�1��G)M�`�%)��Ɣx` �W��E�0�L���V�(������xd�,U"��m�Q�a�C���2�(����>�\7�84�jD�{�s+�o(%�S�������hx�l�=�KJ�1����r"��UO���f"g���7�+�����pڍbXLц�.���i���i5\P���C ���%qZ_�."�6g( �����;��-��`fҠ��ٙ����S�}GSō<W��i���CFk(�i
2��跃�!��F�-���J��V������q=�ƛ�a�c�j��\]U��0I.\����8�B���%�}��v��A*���xw���20������oF�ʌ_���?�_⎐���+�W�n�s)s�e�,�b�nBx6�<��Y[�'�^=�v��O]a�"�S��K5�xz����K<��Ucw֐`r�����Z�ֺff[E&:=LmJ|4����,m�P��5��<�6"���c�[���b�5����58�wmx=�WX����6@K��ntK�y�y4�LL`��Z?.�}J��	w�-��Tm����Q6������}��<J4|1F�e�Gx�� �P���٭�����"|7���~�;����r�I��4�/$�8��S~M��F�(��N��yڡUYL5�b���Y��$*������Rɓ�	;�/�O��i(<L�f�H��6
��Ү�b�e�޴5�,`$9���C�;9@�M9;
�ݘr��o�ˋ�QP��n���2�pF%�ޣ�d�!�2Da�jĄE;��R�R�#��i�ڊd_��I
A��5=L� 4M9B"���U�g-��Fd�2���|P�wþ�*�R��p�ތ30�C��
�Slݺ(k��|�I����A���i�
���s�f�tdoa5S�/��+��VD=j��'z]�ܕ#�ZH�L,T�~�2�V���ϛ�I��B�'��
ԉ>V�L������e�7-v�A�2\Rh;c2������-����Y�|@�x�<�ekU�+դ*&�� ��An��]7�q��^�q����
�{�w����1u�]s:=���5V�l��ߥN7�����v9�<9;�&���hj9.�7�hfdj^�.QN9N(��Vo~a�3z��\�Ԁ���d�w�ۊ+�d��>u���|$��:�eczn��������*���Q�2�ʱ�cT�x0`(���/��)��N=q�3Y����,�8���=�鑀?ml&�s��+�i]�$�v���u^ĢF�� �Ӽ
#�f (�Rv��U�Dg�c�\#)դ���Q�fW2��VfrM��9��� %�+�4zO�	Fej����E;������1�9�ϕ����]�[h��94����0�,��h_��.�B|~ ��\�p�����.E8�}��PU�(�0�F�$C�]��QkQ����"g�z�U�S�w�h�,P2^��訫+�+�F���Q�o��Kp~*�+�#���2\���y� �\y��ŗ`��0��ƹ�W��_�\�4��Ih�l�3����iU�?���kY�\P˅YG�I�P݂���Î�[�f�F,��y�RvU*���	�Ev?5�~{]��j�h>WW��pdr����\�f�m�N�Q�?�����Ǵ$h���BT�I=����q��U�#Mோ,�������Zj�PZ���1p��"�X�	U(L�p(��<�@ù5׻����y����==�hҫ&�3#���y��R2�8  r��B��E��^��{�5]P�5�m`�O����f5�űP&�:b�Nӂ�g��k�#�(�D���{Q�'��]3�o[���mGN<�;��ͻv���Ɵ{�>Vl��%l����l:�������Q�0^�������7��IN��{�]CΪ���U��Ŵ��r�dy���=+�'G�d�)2��@;���t�p�@}��l(c�:��´��Ɔ6�yށ�����G�a�����GV!�̾3��
m�v!��@������&a���ZIXoc�����f�DD� �/\�Y7�d�]�U�4a�����(_p6�����������=[%��;�����)�Aμ�4�!3��e�r�tY� m�B�~<s������/���Ns��o�bjIT�dT��q�ЩK;�����V�g�D��~�:�q��Y?�CE�ns�Ǯ�X }U����<NU*9~��Kz�,H8�9����L�OhV���1���b!���"Y������	ao�ڡ5����p��Re�0������^p���܊�A2Qn3��^އ��'i��
RJc�1љKdY�>Alg��C&]������-<�R�W�\ZW&5��e[3��,��p�݌'�h�s���r9�w�:�&�o[UE4Fc���E?�ZB�l\&2�y�
{���X�TؒF!���D0��zs�iM�i_���\�B�v��q3��J9z��/�*�����������e�yt_}�ɔAQd{��:I�aE϶)���m���kY�go�[R�p�
�v�j��BWow��;�N��W5A����6��V����=!�q��yP���$�o%���A�H������o=���t���? �����U���-J ���X�S�#�S���HK���i6�H�� �&x�*�{K3�X��@9=��� ��_1Y���*\�-���2 +� �b=y�K��F��y��-�dz��J��ޜ����{���uS-�
(�6�}wdf���4�[�ͭ&�"��/�[�Y�3c���k/�����Er�B6U��Q�M���%�?�*���Ne���huJ��5ͪe'�wiJ���ȏ�X,��Was�8/�L̷F��o9����]�0��SJ\�y�����NI�;rk�QJRrE��sb�����ڸ����ÔVֽ֩�/�Ţ��W�`��F��
�.�L[Ӄ%~?�v�UQ���_0J&��~�@M�h�+r�$ZM����  4,�ܧ����y$�����Bb��H�ލ7Y�r����S�S�'f���*3��X�b	�nu;I4w���7ؿ�)��N�u����3^�#��ɈcPXC7�jտf)s2���6#���Hb�%�h�<Y�/͂��5p�U�(�w\a�z�$Eg�*�W4c�`6h��Ґ�p��`�����s���{����>ɌE�E�˾s�t���l2��Pr���ιL,'M�==�G����&�Ε�I��I�ކ�L8�脆P���ۥ���G�_~���@�F���_�綝�r�|1Ȇ�C��Y"{8����.v[`y	�[`�\or�n��hN������ŵ�E��������E<FR��Ϝ�7h'X��\�1�b�3�$�1��C0���Q��̭��x.����'����u�Q�>@��S-'5�$z�&3$M*�[�)�L��#��p�)y�ya3�'�v
���@�W���������II�����	C�-�T�؛޾�侻��L�(|d�|�}Τ�`�<�N]t�j9+��҉=����B��7�s�P���}d/'�B�\
���(�Š�����e�ܪC������C�����9o�UH4	;E\ń<��؄Y!��	79�u7\�̠�d�N�$�ş�>�^�L�G�}M*߸!�󒙲��%��;P�Fj�߱��K�p�ӑ�c���=�y�bA=2���'>Q_�m�#罫l1<����d�XW1+C���꺕79w`��d^����A.��-+ہ��-fr���N%���~��tO!IQ�L��d��M����掌�I4�%|I+�uJ&�5Ec|����F���z4mg���Bj�U�T���jLt�Q���X���W�T�뜷0��_���Ŏ���"GoOt,Z�2�B�
d��:9&��3z���]�;��qJ�|'5O,�������aH
���{�V���?�����L�:�^?T�t�{P�Ck��	Z�J���E|�q�y�7�x�(Q}C�)z��͆���%�"=�b��1�$�����*�)GtPn$�6(�����#��C�����e\��荽DG�^ir�~|p���H���M"�2���Q�=�@�)��Ȟ�AZ���z/֤����Vr��A+~$���bk���Jw�.Vq�ݽ���q���k�3`�|��8�5޺�꽔��'�0ו���y��u��ٗ����Ծ"%������x�9'�`ѵ\k�{c)"pz9�*?9�'�L�L��j��;%�����@4����Ml�/�c�A;�D�M�M&D2��*�e!���$�0G�x.�cԘ�y:��W���WĔ��IGi���a�k��9�T�<U��u)�k|��u�`��4�]��J�6p��]�B���t��H�Xp��inJHJoQ�8{����X����R�ߐI�����Lt��͹in�N���9ý���U��\�WR�1%�yⲮ�q*�W�y�1��H��8ED��Z)��z�p����PZ��^�_�	Uv���[TΔL�-I2�Q�OQGiYY`��{�@��R�7��E����h�ib��&�ˏ����W���k/lc�2z����/��Z�0��w-�>��q�%#g��sA�y0�׭�GkFק�%��'��RћBQƕK롶<\�Ro������&������2#�J<@��i��j~Җm�M�]3�+ܒ��t�f��J���ӎ�-�\����6�r��#�'_��4�`��4�R�.'5Y���A\��I޻'Ц�a/ܹ%q��X{����*�쬆mD�$U�d��_ 6���F����8�w=i�w�1���0�Ac�M9e_#�Q�Ŵ�[�����J�d�*�gS=i *8�ls�qmQ�t���,h��|���xb�M�W&�ȭ�R�ĞBb�M�Ө��%R�)�;���E�h�ybX���.����s���S5o�e�6H����䱓[j 0C�QaG\O�V�ˇ3��Vrd	qW��Ҭ0G)���$Wqb^�kfE��g%ؤT��KN���$Mg��e�?�[g��caa������$��l��H�%;{�35r���I�{��}�ID�("�đD1���yz[h��u4i��zI�*h��8���#����W6�~3I�Nwz�2Q��L	&<K�����T!3��4����NA�/��%|y�� �J�8p�A����$,Q2 y5kdIh�٘kD]�?���>k�Oj� U)74�!kuߜ\Ld��d$��E�� '�+�_����d�>hRה�|���%�j�xa�9v�� ^��X�WU�*�_�DÚU�uo^n�!%��ֈ�y�=�pn�	+$�{눱	=;�,�)R�N�G�_���,G����Q{����$�N��Zߎ�����1v_w�LOV �v���$���`���� 㧀Ķ�R�N]>Ux�X�z:��θ�A)r;O-�O���d2����n���'��!��.$>�Ƥ���9���K��[j���Y���E�l��0�5�O+[\�W�=\�{���L�f��#�DVЧ����hk�_���2�J�#9�H;m��c�X�32�A�CN�|iȫ_��X�c~%$��y����]<�K䭅, ,O���h��6mB���E�CŐK��Y��0��yD��@X��Ҿ���D��������)hV�F��7�(�Vu
3/�q��Ҝ��n<�{Jgv��ft����q�nW:�>���7Ú-��"�����'��7x��G\�3$h�>�kw�}%�Iu�zDCH����8�qsu�����?��&G�8���}\W��`y��)��t�mL�ċ:p�)@6~��$]$���,}D�߲bJ��I�_�B�����G�:���xF��w�D8�摰ջ
?�o�y�=~��ɌC�>�S٥()��֣��ap����Z��!(yQ�g6�����_xî:����BdI���2��-�Q?�?��JQ��Tq��F���o�ͽ�e�,�yM����7���N�P���ԧ0�%+�����= o��-�_,�y9�-�\�En+֗��δk'#��X�����)f�n�+v�mv�Y�x���0�]� m�)�B�v�NC�[Tߖx�H�:~�ZХ�C�5�� �O�~f	���=/D�Y���ɗ*e��j��N��<:�N9�*p�y�C�<�^�X���VC�Oi�`3+��ٵ���gu=.-�k�X������	�����y���B\��S������&S������J d�d�Dt����t��J�&}�nt(L�S��X���n���L�0l��yb`ʈ��Q3R�jt}�3\���r�T���x��XB���D-w��t����bժz4HƚBJ����v��ˠɐ�ڐ��2�'��-v�1-�C��c N�����e�W�v���ՉE��E(���(��߾��g��&𫊽Ya�D-lH[����t����w�gh�A��֊p-1BC�/��NcTӡ���Z��A~r���M��,�?+������s�����7��2��P��@'~{��z�kE� ���3p�I"xӕi�����ݲ�\�UnDE��
ć����ɦ�Q��	K�$މ��'�6�V���@�s��0=�r�~�Gw�=ֵ�M�3�!�'��)GbD����
�;������o`Ry�K�x�?Bɶg���Y�e)s�������]1�*��[$�T�W��CC���ЅPp(3*
	]M���q��e�Q�w:�Kȟ�k<i�-�)��)�H����=H_��?�Y���W�HD�ac٬� ������������R�aC���*#�+¼��gGH�4L�6��x�S
K��AG�<M�2�.EN�k��<�,��j���ۢ�k��p�4�<2��X�c��I�W���tm9l��&���c�7̈́��;��HOuVs�����R�)�'~����ϓ;Id�A0YN��X��Mr��`�-��.9o�Q�0�` �nـ�g"&�\-�=��'��&S��>?���*S6���n�+�ۨ��x��yj��*0���/���[���ýXҔ�J�&:�,	��eH��ma��̱���67����v��8z��`�B��/a���>�yҠ�f�8�{����*yx�VQQ�'f#��#Ac��a�f�Q^yS��O��P�Ry{&đd�{?�J��6���@X[U忡@��������7���U�7��,9�\��3�����"SRp UN?XN�g+��c
6=������x��u?���N	u���"�21 |�����>]�u/��4D�nEݔ��ʴ�ĆW~��NP?�
#����RD@�P�#�볷xʲTK2�į����	t���&a��\�@�섮�v@��/�mTG<�	�M!�39���RN'�ک�O|ŕ�Cj�f\[D`}#)�(���'t�`R3@IQ��݀��<�Ȳ��H���A�E*n�f�WD��}{y�jI쒿T�Ru�`܀Q߹h�Y������=m|)JU,n�tћ(i9�!c�0�uan�<B��v��ǖ��V�o 5����HdP@�����s�Q���#	K�x�e���D(��L��8�u$XoÆ;K��3�H�( $6��Ǉ�4}�OM�.�0���ʎRu���:�QfE����3O]"H�_�/g�wU&ҙ��"Vk*�)ϝK	,p��s����Y��d/bW������Mz�
�9Y-@���l���Jw]�=�+V�$v�=q6K��nϡ��m4���a��G�־�):�VT���#�H4���e�D����!]���RE��t��t�婿���=���Q�Gs�v8����Q��H�x֚�R���n4D�L�Lf�G�~I��Y�}���������S��0��9"׍��*��t�|\��H�.��'�z�E����:���RKQ�9/��ۡ�6s��5dڗ��B?�/ו�jƄut�ͷ� GH�Ϣ&�r��R�]{0'������Z�˺�S���{����B�&�@�vӎ��J��{b�Ɩɮ�d�?�3�JdQ*�9�*�1���]���5��S�k|�`�<��[�|PF�1(�vV���X��V �=�����v��f�L�c��s[.]�
4���$��F��6a�,���/<=����/ 	�ݑ��_�A��Eu��F���N����ϥ��	���R�C�/�r�?Ӷ�w�"
�fп�̃j`Y�����cb�15�L�
-{Ůi��\�J[��𪏺��X��W��b�ᴐ���C��E�����b],�m��C:�'��]XA.��P��95p[f'#����$�'�[v%qD� O��g����)q1q�>�+i�w� �O�&�>�i��/sg:[n���E��wɛ9������s����i " +~S��Q�oʉ!�:��������^�5zIO��!j�	�z�N̓"��%>���|3�p"%O��N�Չ
��u9	�[�dy�41TZ
�IxΌlж��
��b����1�9�X34������� �t_������o�W�7a�0�E\3U�|��CX�Dt4F%Ϟ�j�&{R�So�� ��捤X��pWЂV̺��2�uM����	��+֘)l\�G���o;��	�9��lѼ���P���z&�Fd���`-�����h���i������HG*�#kO
�0���O=s1g/:�~�������;QV�(�$cP�p���A��[��nc�_�[��}·�D��`�Y�y�'/ďjQAd:lD{��q�W���a��yA�:7M�Z���1�L?�BAtѸd_�MZ�;�`T��!¯;�D34�!C�M�"Jn�ΤjC,��;"m�!�(.>���q��x�,s����z��ܿK�Y��珮:�*��R����c�Ua6�ocH��k#��t�:5[Q�	�sdړ^h�]�x<��̴���L�0^.���~�ے-� ��6���*�-�+�7�xW"D�s�����!�ɚX���vO�ؙ�q�`���C��~��U�X�S8n��#X=�W�V�S��פzf���.iUY���72�@�z;̭3D��5��*��W�dM�_�0ߵ�D�a L��������#�ќ�6C��Qg�R�åd(���W%�>�QJ�?��\�j��A�=0<o.H]d4s}��o),z���F�^s�R���j�����������!��e���TG�9>�m�l�{V������s*�đ�?��Jh���6)X����i��z3:F��J��
�:F�f��	/�x�����g�����!��f,�ܨ���"� aM�/]�h�%6c|�r�X������ԋg�O��^���n7r��ڔؠkb�|�[aM�M�+�Y�Ftd?o�N��4A�;1���n�"��:"�9(vj�1�-% ݸ.�~B�f��]a����ء+��^����^�-�א5�I��ߠ�!H��, �Wu���>�"7<UH���y��( �5�g�/���z�m=�7ohe��"�t��?]W9j�v��(�8�����ɓ��W�A�1���!��4�~G����Y����[V-�!_T����T�bN�{�����z��d�D�����nɑ�m;����R�[,���F�FF�Tw+�PT�q�5]p��{>� �� ���EP�-����s�C�#	�RS}K��aXr=�L�@��\{�z�@'�l�|i��ܚ�6�ڧv���X<5pC&�6����D���l�^֢�mCn{k���''b�#����)���$>�5�?��;=���<�rKy��D�h��˝���W0-��.������B��6;R���vChIa����$��X�j�
�g/X+�2�t�������=:/5���)�F�Y� \����XO��+��c�LJ�����;�#8Cҗ�o��U,T_�><�W0��f�S�s�c��|�PNR��M,��E���xG;"@c�J凙�<��NQۧJ��f$6Vä�Og��ǻ^�o9�xeG5뺗�ec�m�+�!����̛,�dN�	�h���\QC��|j<w������nt
wb�m��dgb#���"Pu�!�Z����*z��g��~��@=����M�Z|��4�$t��p��x����A��k��<�E^���0;�����.�����?2��M=u�_�ARFSʸ�HP��/�~�������B7C�H�*Cա��9�
�rN\xm(@C�3g�����rDl?�o�F�m�93j��N� J���v/���ȼǍv�B:L]�d�籣�S���5o���#�*��[�ܵ,)�����};��C�	�������s.������I#�=(e��N*$bP��z'�x�OO��=��3TǸ���zX*\=>�	���Ү�5��ԫ�����\����r<�Y�y��9��&#?�ey��]�D�Z������m�(�wt"�&	� �6S�"00�5��3�+�鰋(��@�I�a�p�؂1l���lfP�d����M�O��^�[�_�����y�$�>%ݳ�ǚ�����v~�)	���O����]m��HW�<����P����4��u� {��̶1AY|]��N�K�2qA�9HN��4����� 3�a��=m*��
_D �e$R���g�w���Q����m��+�_���+"*�ա=3�d���N�D;�Z>,���SYd�	(/���a��=�E0UGg�*%ר����N��B�j�>�/؟�͚<쫜c'$sAVM���R�a�'�.lֈ�1wq1�'�k����p�W.2H�S�tD�-V�/ݭ530�Ef���Н�9v[gi��"��E��n-ïBnML����Z�TS�@$��^�~�{I	vj-�?Px�~��_�c0�ͺ��ó)�M\�Y�*��$��rs���C�r�'8R�F?0S�z#��~�%]�;��8#�Z�Ӈw�^z���"�=<�F��x^��cv	>]�,��=��f������5.�rpXUV�O���g�?��E�/|3���j4�"Ù)���\̫���8�7�(mp�ˑCi��tRt�pJ�~ӕg�b�s�q��v[t�6ŷ��Q.�,5��B^��'�w��6�(�(�3��U��8F��l�c�8:^~�/ON�����a5C�� (��\����ؚ-�ވ�10�������$Jy�`�^Dn[��t%VXXc3��D��B/�y|�0��>���<�X��+�}騊C�05�`=���rR���w�sq�<�w�>��̋Q�܋F���n�t�r���y̍џ�#%cj"�����.�J�9�T�)~R�e��,���u��6fX��ʣ'��%"�T;�v�X.�3>J��;�t�Z�fk��?a����p#�j���$*6�肦7�H��y�c���G��5�|[��}
:����Ě���+��&�#��c��(��\xC<r�8��� ���l(�}1#�����r0�RT?xى���b�͢v���b@��E4���[�����/��9���Y�U0�^/��t�S�=���m���e_�����r��h��ZHԯv����gS�_����]��w�H�E=.�c�a��Ք�Ԓ$����c�\f�-�i6o����n�A;�mZ���}z���@BCZ��j�`������C�AQ@|�<����qB5�����R��뻅�\����^$X����y�8,%�L�D.�>*�(hQuu��[��{�g"�؈��ltYr��~}��U���^w�o�L��/[��t�8�3�@$���k�ݟAN8�a	��h�����G[h��:��(�l^��>*��G�{_���(�ir��o�\��YEv"��"So�
r�*4@7���2i� ����#�%�Ϩt2��$^#�%m��Y~#�<��.���u�%:8�mX&�5� ]��^Y���P�
��$DXm���_
� �@�q��� C�
]-�|�y�������a�#N|��s}��ç��iѓ�m���C)��夿�.FJ�:��v"ݤ�n��;�]��w���W4F��J0r�Pa�|��"ξ��'���O����/>a6�&��u�Im�%1����	�n0�R����i��q.�`�S/���x:��_� {�ُ���S޵�.�A}6����2������"g�km�8�{p�&���W�O�d�1�^���z���l(DA�Wpɹ�X/�s�v���*�g�,�YS�n�y�?�²�Ґ��}�Dl�� 5�K�7!��U�ڋ�������Z��1�<�`��r�ނ�#s>��65~d���q&cŊN�
�"�'�eԮ�3Φ�O�>��IӑF����T�7�N�-x���a��O8�ǡ�ą�ȑ�i~��d	uS}��L�Ԏ/�OR�!�Z��0'C��[N�ɝx�E�!c����or�`Oi��A�����7����S4Z�2����c2�c!@���%�O]�2͵�%]�.��V�P�B���"��v{����������R0u�7H~��L�2�-��-ڐ�}��!E���+��P�d�/y~iT&쾾�Lɲ޴r����Nf��3=�O��:=���!�{���Qb'�T��Q�k���np�Z�E~(��̎L'"�-��8������&V�0���5Gg?z���*��r�vV32�Ht�/ �<X�!*�$Y�����<V��Ci���1z�J���Aѩ]���}NBi^�ɲ�#Ε��ЉRŐ"�sޣ1�4)CD���b�J����G����q���`�p��`SD�7P~�HX)࣯"b���TmσpƋ���[9���>_�E��lt$��0:/R�1+9������/���v�9#u!U�l�nj������2�#mrDe5r�z�VŨ ��1@�/hE�B��N$�����T�Ƶ6>hI�O�Z��`�r�����d�d+�����VI'�����CB����(t���Zg�w�s��3�����b���$r����=���d�F�b2�!����&(.��9��un�ZZ���s���]�+�]Dgf�~�\��Eku�pw���=�׿ ܘ]���eѳ�:¢�c����3�!"X��r����_�6@��[�5�^̈́�&�$e���^Z��K��5I������H�w~:��^���������tBWΌ,�Q��T�|G�G�춀~.��P?u'f$��)�iKqU�X��6d�|˧;�r_@��/h bI�p�߆ƃ�$����Z{[��,]��եЧh���R� d�y�XOq��J١�ă�����@X��j�A|����-t8&Yo_�Qk+�Ͷ=�Kк=�P��dO,E`Z|kYVYd&|tt�.3�<#��\F '����z��ʬ������Zo:Ë~7>���} ��Ju�|6��-�6�l{�
�D:��B��r�X\J`�#�x�^����ݎ1+������P�YI�(�����R�^HH�<��HϦfʗ �������z�v$��ag>���V��ǷkW/�y��sZv��V��˶�����T��G�I�)9�:}�g�Z27_ULB��2\��5�d��%��gd����|�ڃA�O��v��s���X<jg�~�{&����z�*"0��lT��,�d�8
�g��d�G�}�+0�$�^�[ c��*��O5[F����l%��V��'����ߑKE)H��p8�CvݮAp�U|�J�A�Z����),ɒ������v [���c��-0����Ƚ�C��RQU$d,RD#^������]�v=�(��(y���Oi���#o�ٝ����Cn��2r������v赾Bz{���6ĆWRLPERbF��"�d_��
/�]� ��34mbG.�%�S�a�cX� ��,y_DhENS��!�d��w)���@�{*��n����	N����d��)�0���L'r�S{-��<�>���@���<�%d�wv>8�B۲�3���g�� �&�X�:�;@v�s���r~l����M���&��wkrrRt��k�����j9N��9i�׍c���K�y��郲��|\՝c˅P��{*Qڔg��/�or^�?.�[քh���̻r�������_�@��4�=��Wm�ǟu�3���f�#��lS(ьvk�eGsu_3�`����=PkmK.$-�z,�o�m0��0�2Y&��F��&:Xm?�d�S�I@L8DM&
����%f<����*��Y�G�by/�~�J�l���l8�4�QHBxމ�i�/�P<�8�;�^���DN�*Я("o�VKC?A�Z�g��#l�5�N��o�_��`e\g�+HM���P=E�'p����[����j_cs���($
S�ƄSt�&�ݝ�W��}q[T,�`7��U�s����Q�T+еjb��
�}y��ʃ���Qԇ⿅G�|��-m'���0����G�Y�l��G�ى������b;i�.�RQ'G�O��X?��i� �p�U����&�N?��N3��Jg���'")F�2���?�_��-|ibx���u;���(p��y/��S�1���]=Dz̖'.̘e�y��ٶ�����;ۆ>h�[�����Ƚ:M���~������k4�tY��?�N�쨨*By�+=��T,���ĸN��I���P��5eJn���h�+j�H<RF�V��A�u4?����\�`�Y��1�����
���CCh!��(�Mm_�c|������E��
HF��D�RHi^���M�"[�P�9}g7�G;�� RAOH?o2:��Yڸ���N�6�b�<h�Y����G�k���ff�&;����"Ӯ^b�O�zX\���
���'՛K`�&�[��C6��Y�@�.�[��*�E�LSh���\�rS�9���cv�E6�k�:�ק�F�,�B.;}�������R�H�p�����|�U8�\���d묦7z�q6��	�g�������E]GY[�2�����Ά�� :�B
�)��.l�F��g��j�~�sJ�XM��ŁOB��ىDP��(�AY��/ZXj	��Y��6I�WW��Q�	�����Wd���LoQrY�8[���yɖLw�,�Kd���T jtݕ����4�F�����n�_���O��>C����&�W�Rt�"�:8`�a�\Kkv��7B��P�,< "�/�-���=�ۍ��jR�dEp�9R�GQy���?�����vإ����h�X��+��,�x!���]
�ďRu�@� VŶ7@�RXE�=��n �m�ܙ��σ<�/߃�jґ�hPH���=t���N+<n\����2�Ga�7T�?u�� �椕����a7�9�j+�t�	�s�ЈV|
�*�E�$a����V�S��,���E��`͈�Q�ɔ�m�
���1K�@�3j���9+����1�2�Mf9ǿұL�p��<����+���r�!�e�m���HpXs��߿J�܋�wޭO���kS���?S�*�B��^w)T"ڷ���%������$�G�����~�165z��P�!�dڽ�e5}�:�����I�[��ȣ��`� ���.�-C�:t�pZ*BV�-��B��ܐ��v����H��¨;�D�=��+�/k(6=`��,96 ��`x�`
�~������m�K~��nK���غerp�;��J���L��b�6$Ri/Ӳ������!��<k���7 ���	I�J0��8�q�0��5��OX�sж�P�E���qD������7�&Pex���@��A]�[�0���O�����c�[T�k�?d������%I`�ǄÂn���zdX���״��_� �{]�-U"�Yڰ����1���>&���4�O>H�*���sKF���A	;�P�y޲�
,���V��\T�0Y&�A�KE2�-���x#t9�hx�_p�����l��7�Zb2ly.`e��-m�.�@����^���l���'#�W������G�ۙ�$椚+D��dE��n����g��G���L�Y�qAȕ��U/�c�������)���d ��a�&5�C�i�~sH,i��(3a5�����5��d	�u)���?����N�C.�/��,�N�z�nP"��<��\�G��̫�s��Z�j��(�YL�	ƍ*�F."���SƘ|8�i�U���N�X���D(L�pG��T��5ȌE�ur��z�S����>Z3>}8�S�_��K�;�׾G'g	���/�"��mo8;�͙`�r���ma� ^��B��ݞ�T��E=�{��zQ�5���HC�.�{po������θb�=�a�<"��h�Ԯ�,��w\!-.�jn��a�β�B��M����^�>�C�0*��T����.�:�/̜j9���T��J����<��N��q,{�p]ld7M�DR����@�Rj��P�ŵ�pd!0���Aґ@(�/*4�.��?�8��J�D.d�v2O2OP���ُ1�U���Ben�L�鮫��9���]���?���B��S�	f��:�N4���@ʁ+���y]:?���h�Bξ"-��ͩ~f�P�,�M�BW���{���NM�y�xI�����|a�F1m��y7��/Ok�;X�E%o�'��� $��[K�n���+Ȳ��0�2�(�\3�6Ƭb�U1�f�]�	E�ց;�yº� m�w5LR�a���t��M��,�;��/�{biG�}��q��R�Q���o���|V�8����[�Q�j�������d�J�a���G@�]�,��Vf7�����A�zG�ȿ+y�^a�qb��m&�a���.��K���=c��� ��ҹ,���i���G���+s��?�'N���j4��Я
 ���Dh�]=Zw(d���ؿ�U��!а1������Zu^#���7}�a� �����IA���΋>\�Y�ɢJ�Y�]0SF��G�H�$ Fh�|܊i���d�d�g�3��M��뵋e��H�|Qv��/��{_�oI����j���
��ereźR�n9�"o̓Y����eK��	Ey�������Φ��� �H��32�����#�|f���\����4C8��Q6Vb�f�C����
)kǟ��CF@�+�<a�\׺�4h�ͨ5��cر��lr�G],�B#MW�Z���+��7��9#���V[',��9V%Y�I�{jt�Qp�L�UTzCʞUﴬA�R�PQ1�7�sތ����0�!� t�Ip��إ���,��{�*�EŬ2�X�F:
'fI����z097�7ȋ�-�H)�8��H�3܅�&��Z
��Z*�#jA}U���v(��r��K4Ŕ�S/� ���;���P�{�V�����+����+��r\� U���>g�9J�H#P�j��|sEQF�=P#A��V9
�3б�W�iojM짴��π�m�^Z��S)��a{��b$�M�xV���NH��g/��T�R�L�$l��n'^U����z���Z��}H�#Oe�	�K�u�W�f�#�N��]Z�'��
X4a��a�0���Ÿ�����l�=��0�5d=]����)��6-��,�(���0��
m��co��@��;�*�r���>l���m1��� ��?��;�~j}�Z��Z��L[�͎y'��R}0��/�ȥ�z�g���Y���%�l��˾|'<�N=j��z)����E{ݢ�~bB	��`�(�����Ws���I՝�w��'"]$wc&'����HV"T�s���mg�> ~�΀�T����:R�g
���X�(�LA�c{�A͑YUҜA]Q�Co��?
8t���3_rvx�ٶwI���D9����Q�D�ާ ��e�?j���3�zA�Ub6/��ᖗ��4�wN�Z8�$C��ff��`�Y�w���,�a����{q���l��ڧ�; Z�����H�̒���%=;D^д ��vͭ8���%��1s}҂�(Xgr�R)PF�V���lF�@��|�鶭r�L�"��ȁ��L��"����Iw�i:^�M�~[~z��Ό��vL	�5B�s���������K`Tn���)�B���9�l�c�����N��c��.�&�C��t�;ʰ����0�͘�	0��ϴ�.o�it��O�C�U<s�0E��p���`�:%����~�l��/�w�3n�g1	�9Zf����g��*`	t���`��ϵY�"��9Y.��j�*d�V�)"53(���f�hfG�؁�رGR��z�M!�@�2�Դ2{.kz��D$d��m�[�X���<��\'��[ш5Е?�IG��H�M�R��c���~@51en	�g�6N&�0J8�K �G�\�EK'�8�SxD�AGA~�7P��<!�:�PA\O��/�N,�>�jݴ�K�VZ#"�X����5�P�ՌÀz�X[O����x�@��F�]��`Q���}��L�e=���eBO�̔7����t$�țݬ?!�$�:�KS���)SL���'��yN�h� r��nP@��r^���L"].��ΈQ�
|��jp�8;ü7q�ޛ�i��F�=I��"�y��Ǩy1N���?/ac�@M=e�:�pn��d�j��a�9Ʒ���'�2��ы�Edb��hb?Ġ^��>@@�)��t�i���@HFk���i�1q��ș}^ck�$ң~k�1���(�cz�6CV����n8|W��BZ�9@%���NI���"��Og����g�(��Ѝ|si���A�?G��5j7r�����`�3M�ԁ�A�9�V_����.o������:��Dp��=>)��o �w;\!��Z��1�����:TD
�P�N�[�M����dv���;���9�)%�yƌQ�MJ��*G�7�T���J��F��Y�v�G&��~�>�.~
T*��r��@��>0"y��z�,��x�_���@'n>����X�~xd�7�l�-�s�w�,��u��RV6@|��d�̻�ĎI���n�$��=s���5h�?�ar6$���V���I9txρ�i�k���,��2�{�/�ۢ�=M�{Bnb�,J�'��5�X�p�]�S5��%�?g-Qk��+�0NPb�b3�h��
��m�KWV����������z,ʟ��yH(Z �2���Cm�.�� e�R4��Ґ?����A�ٽ��FsӇ�Q��q4�u*�)p�$W�ߝ[�倰��Z�S�&��
�9��0����/���p��5C�g�,C4k!����(�/�/���I��+s3�"�\��I�6�X��[�~<l͢�rR%֨��IG�k�D5�X��ʩ��$�]��U�b�������f�����B�J�J�\`QD�e~VtS){�#"F��{̂r����,�^Y@
�|�u�W�B�����}���%����߈e���d�ũ��S ��sjA�/	q����%�#���b�K�#����þ­��գ��K����׼���_C���JK4��!4�rv.�٫)�s��Yvp'Σ14��P0��I�aI
%�~�N�EN�����lz���k���((���}�X'.�U�p�����eԊO�yQc�hlA㳃_c͢���Q��>V!K��*����F�XvĚ��f�ѻU.{�h�A�(>`r��
�����oc%O"r�#���.�����*S*1�F���$�u'$2��1s�3�hc/I�����)�/�Yw\���o?-}B����&6_!�J��t����;�$�L���rnp�	[e��`�/@o#H�ް��`�8�y�Vsͽ��<�볩:�D��~K1��;F.d�A��[0�*aEA��U�r�ai�N��D�I�&�&��ۖwZ��%��>�\���D�	��<
�,��c���L@H��a�2�Gi�_ z� xÏ�a���a� m��5�M{c,�%b�:H	M��ji*J��0��ex�4P& xf%ub��WF�R$F�(1(�3�j�b�TyƯ��keR0­HM)�N���q+���
����W�r��V��ߐ�
���X<��݌H�<Z0?߇�j�+A1�6�sq<b���9%�H��o���Bu�y�����Y������:�ݐ�Sr�O59^ݵ�8{��\(bE5�G��rjw�[C�\a#Q�c;�䄎��6 #�8�9�e�?"����`$r$�(��c�J|ЇԻ�	d,�,p��h��v1J�ڰ��c��K���W�+s���T�?b�jw���������>��bh������t��Tl�H�h�x�^k�mU#.��ͽ�[IϩҰV��
V[EM���R��e}]%�P���2����n;@�t9�n|e��T{/��!q3�bk���=QrV;��C�t#�����Z"�>Eg~<��cnB9Z�<<���M(:���Ciڇ8d�"�xWͮ���/σ?ݪp�A����pl�U�g&d���ר�4��9�87D��^��Q�1�H23Q&�cźo_G.ou���Hd}+�9��azc-����R���a�rߗ�!u>+��\9�&��(W�����`�V���nX���"�$Ϳ�-���w���-�b�+u�@�Q!8N�VU�_O�YGdt�TCԑY�LL a�Ps%����o{D�찍� Oe59���{Q��ۉ�.���Wd��t�Lf��/��+��{����f�����D 	8�^� ��%,������Q+Z 8�X��0Xk[���gA�M��\�='#� g�?��ԊF�����h8Cehf4�z�pDpv�L�zFVhS�c�v<#U������1:��$7�<�8��Q瓽o�ak_'m��4�G��M+����m� ���:�����l��+T�LTm�u��vޛ�Klt)��y�V��2,��-��xj�H���;_k�Gn�s�=�
�_��H������.�D͝�$�y���>W�ۜM��#iE9To�(K쯈��]Q��Yax�:kkڣy��-��,���yʠ@���/�Ƕ�-s����̂Ee�����muZ�S�u������/ri�פ�WN�l"�jw�ĚH�_Q�%��&w�1)�͹9P$n� ��C�'8��7#�o[���p�E��s�0xM-�"hϭ]z9t�\�s� ]N�8Aݬ5�hĒ��?�w�b��)���l���X�)�����2�Kgb7�L��ڛX!c�v &�!�����90UC�V,|�fB��b�4��wlv����CI�Ѣ�nuȗ�B�x-:#ƞ�]���z|鿵����ʘS���Ew����A��q�{-Mo������-���AJ��~^�Z��Խ<��fY�v᥷A�Χ͙��:f�\)�ӧI�>=�{�h���VK�W�^��f��ÿ�X��Y���,���P�'hYY�a-N1N�\6 ��ML:r2��ܜ��������@鿅AL�I\��rw�v��#�#������6��%m���5������Q��	<`�Gו��E@3p̅�U_�ʙ/.���3X����nܲ��H�9��@3����{���No
���]��j�4����Cߌ��D@��Hn�m;N��g\���w�Z�1.{�����5� �;E�f�%hHL��wS��4�٧������[�'�J���D�][B=l�K� O��v�z� t`]d�i��ۓB�-9�c�Y>�v#����x,j��\�Lz�6����!-����9t�0�O�i�O5�����q1_o����*kC$Ν#�7��q%郄�K�����K��AXw�'�&kE��A��o/&��N��'�U�6�)�g��FR�hq{fV�(R�{�x�x��N�Y
���Ӗ-I�6��P�H�Y��,���_�=Pu�� �@���~,�|Y��9	�:ξz�Nl3�.�.���E���{Y[��<8�S�Ģ+����@���4�%��|����� @���
��Ȥ����M�r~
����'��)��FlL��+�0����͔��|+@D5�#���vc��qo�S�!F)-SEξ2���ߚ$���7��l����4�g­����2�Tf�Tc3M�A$|Fs��y�'�7�5fD����͜��<���b���~:���")�����B&
Vo�f�)�}Y64�WUc.窜��1�=�Uc=��M��"'�E�;�I�h#qX��M0�"+84��ja悭��l{�>&�GQ5�R����y�jA��J�R+ǳ�*hz�09y���~��˱�`����Yk���y&:��[� �$I%��R8P���o���+�����eOh�ꭘe/�g>�L-+�v٘S��M��(�R���T����p.a,��g��yՉ軐*�J\�v�Y�]�m3��e�-ER���u�W����}��������1lf�f����~�1k蜁S�ȕ<�g^X��+3��Yd�8u��J\�.~ϋ����DM�,b9$����J����&����̩U��f�x[p30}���8]_t}�SqO���ɑ&�������>��ż�s�*1�f�{lIB<c��A�T�O�b(�Uڇ~�V���?./Z`W*���� B��?2g=�"� �j1���L��L�(�!��������͸�o�(zn�R�_�0�gR�fUY���|�[��DB;���!����6[� ���[�n[�j��0d� �<�)x/Qa0 ��!ߔ�8�������հ���%�k&���������3}��v���Jp��iZ��',Y@��y�<�|л�lR���Vg��j�^?��2JIr mv}��ޕK�yv/�l:���9{!5j��k����բ GgV�n�c��0#�+�����/t��J���b��lScM�ԕ _�/!`R-zg�l�:Ԩ�>�j���pѳ�řF�U��P"�aU�W @q�����D�»�jZ8-Q(X��T��*� �xm�_f����^8�u��2_]�g�8z�����.�����ɻ�i���o m��?�B���n/����SP �	�z�b`�0g#��X��a!��ذ&}w'�-E��KD`��m�%�h�J�Cm1�q��Jh�0]�$/�/�����ņY�5`���Pc��U^<0w	��Qi��l�C:��JJ�ގL�f����L?=⛣"D ��0@ �V����Tk�pPc	� (�*?��>���;5�~|���H���"�vX�}݂R���+J��W^.�}8+	ز�l����oW�ctx,Hi��@-g����@�[���P�cK�XOQ��U�H�kn���mZi�.߬g8��wl��P�p��yX��.�*��&u�Uw�n�XZ+����|�5��bBڳ��y�}���֞�-���<0T��D|�E�y�U��������h˭E�y��d�Qa�A�ι�a_`��|X�����?�3�� ���'���Ѫ�F����@bdʌ��1�?����!(p	��|�g�mY�r���C7��{2_�!\�o�u������tdQk�"��Ӎ�FS������$�R��xg�Fh��ʃ��m�ҿa��z' �٩���1�Y�0U"��BVb��h��[K��g0�Q+�~��؉���a�C���?�U������"G����ėU{�)à^]�Y�tJ�:�bI!�d��nz��W���� g�b-D4xD��]�A�-y��*0=</͘\�]c�!��N1���x���"�l�T�`6L��Fuf�A����I��Q�Λ���
����7C!Χ�A�cV.��>g����HY� ��*�\q,Cuw,?���L�2�g���2
F\��&,#��X�s+	���{}s	˲u�p&υ{�e�+}@����?�﷨Nu��x�m�;�?�~h�$M��(�\&�����Δ���+����h����LTwv�\� ���
{��q���vd!
́��-�P��U��f�>`����-�{�e���478�����_JÝ�v�}k�O�w!�u>���+=�~igk������L��APN��m��?XI8�(��;�m=�I���w�B��@Y�ď�&��>��M�.��(d0�>�#�.s�E�U��&��Uk���jzSY>=�?��bcϻnT�r�i�A�U��QQF����@ZП!IZU��U�A��)ST U�]<����/��em��)�|���,�y��nf����n"����v
�1T"�q.���$ J�����5ʙ7�$�m-q0p��<X�����o����3��"�[�L@�%���Tu��E�&����D����i��L���v���U��0��yL������ڊi]�}T��6#Fu�JZ-ypK��y�^ګ���{��E� ����Y�Ζ�E�$�dh��W��*�a�XLYn\�l���D8{K���.U�����9UH�%bfں��o#���Z+��>��%F�ǰi�u2r�{�(?8�¢i�*Ob����D-D���!�osY+>|�ݎ�5��s�\����>�Fu��PPN6�fU�Y�[��Y�h��;�:p�~:���8Uλ�[DW�����L2��{��.Y�=�!;�R΍%��i�s=<M�\���%�H�,{;49	d��E��P�@������K���u[al{yzo�gkc_ ٩T�-��b��[╾���	��(16�7K�P�U���z����)��t|Ĳ�&�^-�p�� *���[�c��>�}���~y_Ļ�?*v�}A¢�����2��4b��fq���znC�
@�z�Q��B�0��L=�Z-Lrc����u�w�\��9Nx����C׶�]�(B�=U$K�F���nr1�|@fޚ��>�k(S�Da���b��h�ZxU�K(���^�w�ƥ���Qp3���S�:I�?�2�,䭝w��hp�h��[�,�v�ir;��a���������/�N�k?_� ��70%�E�?��KP>U>���VbBL,�`��������j�{Ϊ?/9�ﺅ��.-�X�rCܥ"���ۍ���1�ڞO<@���,*���$+���tb�`(e�yӧ�Af��������3nspQ�g{f�m�c�F~A�Ƶ�N8���,���'])����7�j6;'F����C�Jq)�:V|T��-�* �ZCZ����ɯ�h��C�nk�t��5v����È�슆7��(x g�OKf� ��X�R:���ɡɝ�Ct�0�+Og�T��+�k���#_�6��P�FC,��>�8#a���-�lI��.˘���>��+�z�V�d���S�!WO�s���a��"�z�I(��w�ۼ����M��^K�m ���6��`JR��W\��ۜu���v�5/d����-Aߡ��H�;"��u�ޭS�f�E�4YX������.��5J��S��s�#��>,�%��HQ��Z��_@��u�}�{ G�ݵؤ5��hM$�^�g{,趁c} ���텧>M��5Y9E�HܝݴRh���iVF��n�K5&��M�����2�O�d�~)=��i�X��(`���&�<큞�0�=�����Ɉ[B#{�Z���C�#T�]�p���-��K8�i��x�LGݰ���Xh�t��`N�8�F��u�%����9E7Q�^�J:+d��G��I�*�o9o��_ ��v��Q��M_����Z�3�[ſ֌��>}z���"዗0�.���?�|�OG�S��@�-<�M�f��@%�C=u�K�r9��wm;���DyB?�:g���l�{��+�{����(�S���ה��9�n��15��B�;�qK��
�r��Cq�2^"6D����,�՚�-CB���j*@}L�Ao�Y(	��nl!(� ��9�7�4|�G͹P556muڲ]/��%�̣�cz����5;�*�fP�pI;��˃�	��-�O�ݧ�����Ǝm�)���g�P/��J|�"ࠏ �ׄ�z��L�"��Y~m�������j��{M
��EL�_��Y&�bDI�ד�ř7�3�w��Q����7��'��Y8�c��P�'�k��b�}�=m$3��ٞ�����ܐ��\N�׾K��I�}����t��cMl�U� JV S\c�}R^o��A���b��,�8�r�4�떖�����n��zI#�ʡ�[�#�+ ���O��a\\lQ(�v�{��a��L�*�%��,i������s�5�O�nQT�fAQ���a!&{��;>	�C�������ދ}lƫ��O��iP��av���h��`⛹�"�9ȹ~Q�.߻lU������`_:Մ�A��&��1}�j:�j[v�4)�1���ݜ��'�#��a[°x ʱDl��P���3����n�xf_H���Z(�^|��Tp�h.�e�n���%��<ؕ�_��hg"��L�4[���o.��΢2�u�2w��~�K�Y���WRW�;CE��R*Pr�T����S���<|��U�-�~G�w�S~�/��=�O�������0��Uv���Ђ�c�5�.����=�L�_�k E����4p�fĈs�X jcA"\��v10���&%���-��(_;#��h?x��뎠�2�QY�i��e��3�Wf��,��;���yÛ������ԅyK`N��bϔ�,�Dd�����+�b�[�����_�uw�(t��1[F`������ O��vwp7��񘢠K�?0[�a��]�[u)K���~��^����`�ZN��|3��|�u�%���fp��4�{G�D���K;u��|J8-L�P1�(r��|�>�{�T�j�����	A��NE�8NP�����="�k�M��>��Q+��'�a V���j&î̝�
��%�<��wZz���*�?̪?�e�ۗoViռ �Lp'?n�{  �#�����u)q�Z	0x�P�#�/y0�f��{J?������簜$��8Ї��8��5O,�i+�+��\�|�$}�V���ل�r�/Q�&%�o�w�)�"����cVm�k���"5��Ld�& C�B��������nx�w �beV�f́���H��i��fg����P�g>Z^O˳Ȇ�kv�x���	CU�g�Ӆ�:"$�`zT��6ȎLD����0��^8g�`y=�5ߜ�K�;7�z��h��Ic��q��{��:���=֒����V2E:�Xk ����w$�c�����d��f81e��{_l��á��"��?��U�he@�>[��F����{���)���wE����^@������ZY�;Fl�o��]Es��2ہ�d��*������Tz�.!���W��i;�Ti:%���1�d���U�!w3S[ں+��Է>"���7��ς��x�#�:m�<�b��b��}?��l&k��<}u)����|S�i���9RluS��Un�IL��V:�O=7�.��ꓭ5�c������Ę���/H����G�`��������߁���kL���a�8r���֓^oabj�$��n��C��	k�d����vl��?"RG�_�2ӑV�K��&�D8����Mє�cf���ND�4P Z�0�&L����D
l�8T&l�����3Q��<���ZP��K�vk�Z|j�h�ޯA޽��gn�Iji(	ͻ��P?o>�n�	�$��:]��-q�T4�Ǝz��$�yC2��6�"�� �(��P�4 ջT��閅5z���s������2v��jB�Ԣ��Ŵҫ�j���uO��pU
g���L��y�)����Є�H�-���2�g�-�X�#��tYF>�I�hb}
�H�kz�E:S��g(���8��d��ѡ�n��}-ȶ��q�D�.oOu�I�<G:�[��5����W	0��MJ�[i��O
ab�h�Z���x/�㶭�k���+Ͷ��oB#n݈~䢗�w�R42�9Jl-6��I��1���.22iG�s=�q�}%�����S2��T"�H�;��;�Y.y��)3av\�w]=DŻ1��/��@�$��(�*0�v��c��7�.�v��ÿe`�N�ԜT�\5P{�)��{�Yk��z(gUU5+��}0j5n�����b�6��E:1��~��[yr�u�7&m�Y���0x�z^��8���&{�S��K��r�f'�\�j� H��-!Ɣ�έ��V%p��`�]����'��)V=� ��ɥ�<�PE�k�N�k�c��5�EꝦ���c�iٺ��uY��>'�Z�g9�twOp���!d�iy_·�\�hw�Suyۼ�����y�G�\��aߌ��'"�
3� �6�=�HR ghN� )��˧�����b�M�fK��V\�]����7�:�C���z�� ��(t!��x���ǛP��?�x�&/�ϯU|�~���l^m�E��ŞK;R�+�Z���������w���Yx��t�t �E��l,i��-�zU?� ��󼆕�}8���8��Y��(�LC_V�w�Kg�*�ڲ 2:�5���^ڇ5��\�%f������K�2�B����`Ҙ�r�XY���]�c�?����˟���Q�<����m#�U�6s��������z��ҽ7��-�6�F�H��2*��P����
�J�V/,�S�(O��_�)�1Ҿ�N]ķ��
��r6\\���Y����,,�i�ϼ%16.�.���k�F��[�� �\����[x~ݩh̝�a�A�;�-;4@0�}�P
,~�p�E2����'|��SP��-�,m�;k��Oh�R�܇�����Tl��zf/$�J��|������>2J]Y5�s���oV���qk{gډ���8�~��eDb��N��)����)�s@���16!��)DlĬ��4p��oK��6%4j5iljqfp��3�ɍ�X�،[��F�p!���
���~�8��]]Ј�u��+G9%���q�r��$��0���"�
8��ɰ ���7�P �޴�;�~^�e[��㦳XpR<�CWi;���:S6�rbz������m��5�X�Ω9��i|��$�HpY����z/C����RT������$�EҢ�W��!���co���ҕ�5�z�'���}*>N�R{a(�5M�����W9�����v#��ד�Aԭd`��PN�W/-!y���ޞ� rd�ǧ����,���Q��Y�'V�k߉�9u�M������p|B �8�gR���i8g����/��(�P�����F%�^�M^�o%���M!�v���.P�'4��hE˓��q>��Za�!zӥ�P�N$A�ڀ��@f�-�Ʋ�}S��j������.l
el���d��0���%И��b~^�T8�G��G�z �o�P@���g��K�.����o]p�=*sF�N��L����bN��(N�1}���ݻ �5t���G2��em<&�=\�N~-��8�λ/yK.�1������ª��6�\
{Z��	@��k���-�)�X�[r�y�� <�R��x��MA���6�A��K>� /`�Ys�E!+8����x�߉F��5|�CY�\��":�D�����Zb��xa)��SjKn��� ��
�<-בɗ��.x��[ɮ%���D��Ơ��;����}/{A���|��Ҽ����Kng���a��r��a�2���ݟ�G�lB��6ɞg���S7Y�YL ��p�l�k�@��{mS�d���� E���k�z_$ j��O�T��T�
��l����x"��ESD ���>l���s�N�1́��`�6*~wO��p�y�˹�R�`S'�nicL�\��x2+3&��������q�ʡ%��>��n��#9V0���GM��L��Y��-ı�w@�	8�K�~!��C�E��&b�UL�6
��b���a[�rhH�*d�o���rr�S05�nsa�\�!�g%$��]N�Ȗ�͎M�Xo�:
:�P��t:lB^���#r�ɕgz-p��m����Jd�/'=���4���c;�#�٠Ex	$|���4�]���(��U�Cu.�K( |clmtى ���=���	�s��,IH�R�·ᒴ������ ��8�W4]�|�1��C��{>�cJ��F��9\lHo��r-ȟ8(k�s��g��.����q�{au�����b������w|�A!���W��@H%��n��[@��ϖ%���WA.�AŠ��n\�[�,y譫���,O��?+X�3ɖ��XOߒ��-�f�'C��'��#���ݝ�kL�}_4lũ}�o��UȀʥZQf_��E�O�z��4���sP�aЇ�� �ʑ���Tg�V���k���o=k�=lF�g����{���n��N'�������_7R�2������ծ �c���6s����s��i����z�`��r���YV�[���7�z���k� �\���w�MT�s��a�P�}��Y�M�&%N��88���k��w�'�%��u=	��1��cd@t`[a7 rw��}%y�%��l�ϽE)���e�0�!�{0\x7�@��u���}n�z�<��+)�2���h:�y�[�@�{'���q�2x~;�PR�T"q�K	-�6o��3o�ҳ6�[r��{w�u!�w���[cN;����O3Q���q7�U�S҅f����PN:t���
_����-�#���:Xh�\"m_j�.��ތ���
�=��W�)�]^�x^6K@�% ����v��!P[1����`�Z1)I�i�o5x4�FM��t����z~�i�6U"�P{�rY(,&��l�j5'�Adɂ��;���+e�U�܈2s#t�����{=��`Y)�����?�n*2�5J��V�8�J*���N'�j�O?ҳD��'�Bl����9X)~e��6.��4���6���Y3�tɈƤ��U��Z�>��	�65�e�ӑl޹�m�AJe�0�8��}��0򡰓YOm�Y�'�H��]��O�xՒ+]lJ�]Ӊ��Y�3H��R\ϸgF@����"3���B(L���Ro!P����GX���	��o�~��㵺�\�8P�C�������#ľvٚ
܂Eo�t!��������(��
���x��ע	�h�ݷ9��Qp]�J/~r��X��4ҿ�X�3w]+&�$�{�4����_V��j��}��t?X>��K����|4%W�MG/���
M�Grr����j]�؃�|��iF4'/L8]��MM�ۏ�D��E_�Ą�b!�[CPt�=��X�X�46Y�0��d�����dz�A��}.�{�00������v�;tq�f�����'�j2���"��:oV��:;�-�e��Guy��4�ɫ[$��4N�!��R��7s�$��>	� T�o��.�� �в�������"i=�2���s|�4��!@g�8��>
�J�:w��T@[���|\y~ y)���i䀈8�$�����3:}�9Y:I�̄�!�G�_��0���!��wX�����n����Y�-��pJEktpk/��t9]*i�|�\! a1O�O[vՈ�9�%H��`����2��@�A���t���}T�;�:��'�ؠP�Y|Ӑ���.:�������D`��m���9:����{�G��nWq#Fr�>5�8Nï�s��;�����HkjIVP�W��Zz�mh��m-�~A��9�7`�g$�"(����{�
��+u4�
9~�������U�@�8����J�f�x��w3��c0h*�͒��o�(�YZQ�<�ݸ��@�g�!AW����������蛷<mZ=����ey�������'�$ ئ�+�eЁX�$@�>�/Ж��n�i*��y�!P��[���3�`�	O+�	���o[��nX�3���D���(�0�F��N��0������Okޣ�0�?��r�a4������&�
�(c�?��,�����{ѡ��i���%�+�b�-���[Q�*	N�/!��آ��'1��17�����O<Ú�xV@�[���Cr'��P��k���{X*C�h�.@S��@[�pg���:K58��R5-h˘F�k>����H`/�6H+��O���~���-��F�e��Jt�D̽���~�l�U�tD[�E�����w�r
���:2=ա}��$�pۦ[G��%��ݖ�zXi��l)�sl�����?f)�O�=��9z:�'�R]������!Yשu_<q���*��s8�P��E�0p�����Y����=�[�[a��Y�6_71��~��o����ػS�l�w���"3EwLE���A}ځ��Us�2|%�pk*���4�e����Q��I����c�����s��AB��;a8���k�"��r��g����O�>�4K���qwd�>��JS����oBJc��?e�"��O��=�	�F�-�2�D�y_��IY��feB��nqJ]-�w�'AIDm���*�e��,�*�֡<`i�h�����r",�;'eD�T� �E$��P2��8Lg���t�=���A_��{r:`&�������d4��wcKF��Z�� �ol��9oX�8�@����
�|ɴ����.��;,>n��2*��9��}6k�9��{}L7H��%�[�k��ٕ��Et��ύ�	�t�A��/��r,< Ϣ����,�Қ�#��i�!�T���{){�*�l!�4���%�V�PJ�
��y󪳽�9Q�'q����د�& �u6G�d�ϜL�[Lz�jy�1���j�>���Ub���zO�S�����1��b��GT�����6j������}K�~�䲟����W��%gn��O+K)e��|����[p���������!�2\lF��xx
���ˈh��]��|54�x���O׈�a&c
~�'�tƥW�R�"�fS��	<B�a�M�b�;]Lp�G^�t�/)��
cpY�����,U�Ǆ�"�3�*�W]��Y�S�����pa@�ͬ4�����aC\ǯ垯�M>�h����:_��+�r�T��AK��Ɯ%mR|��ɧ[TzۄQ<:	�T��wq��墡�����	ڿQ���g�#�I�U�Ñ�	���oߐ6r�r��6j�*��~.�H�qc�����{�����y�R[-�H;&��A������]%�S���\S����¾S��$)��72�=�?�Zi�0��)��2��@�M���DQ��-'>'�V<&���5�Uz;u�&���<DH#��'�r�S���[�z^)�x�lv5&JL������ߏ�]w�XO�ۥ1����Z�Z��f�6:���j4�_�)bN�rƿ]���r9f�"Ο�`�tI�������n�O�/��c�cU��c���a�O�_��T�����U�4��9P^�� 8M\�t��y��猶�I�_��-�%�Ӛl�Q�	X�n��"kFX�����`�{8�;�:0>^���laoZ����^w:@n9'��]z���O��]Z��b��I���}1O[�}�����}��"��+�_e0�Tl�#|pFݶm�fA���YDD��Sܙ�Ha��D���X?�	�S�>0u��Wh�C�c_���M]�>���*�n�uJ-3��v�#��Ӣ%��d���\�ԅNYA�&��-���w���K�֪�U��q�[Z�
O�|g񏃿�#���͆� ��ӷjeӊB+�X����H�=��@�����z��p*�����I�Ƴ���e���l9c�c�k�?���l_��{x���f�ͻc?fu����^��^W��K4J�c�?��W�4��L��F����a�����*��ʂ� ^W��R��H����R2���'�pK���ؠ]5i�B`�T@����{5VՉ2��s�3���j��jlф�pp�݊9�� �5�;�m�:�/N����b�/���*�r�&��uYnCLR��t�R��׼�˟�ȧ0��X��3`��ݥ�]go��3î1��x��i�����SS3�A���ay$P�J�(���Y!"��C4Ar�����jI�*��������G�����i.�
�?i��%���/Z,�Cb'qլ�`�W~��l��~����׸�M�~��2�D�C�K����|�#��x�ےU��+�#ZVKOb��)#E�ޭy��Pć<څ_#�Gr��D'�T����O+�:K]�i<�$���.�-�� �U����ٔ`l	;����V�}�did�f��W;���=	]R�{�`bu�{�H39b�ǚfǯP���y������m����0w̽;X˜� .���U���nMl1�JZI�`��+�O��×s�c�6
����(��Uͺ%��a�l�_x���y?�@�����x�H�1:k�H�N4���+v��x�I��)���YoF�r����U�� ;��G\=��6qG/n�Kw�e�����/����a��sS��?/b1ФBo�Wƈ���KV�X��XT���n.�_L���/^�vS�Sԓ�����Atc��gB� ������4U�u�Y��oytv[a�EM~���&�hK"��i�P�ޞeu�F�a��ۤ�4&�j6��yh������ϯq@�7|���B�1:�BI��{�Щ�)
��o�\h(69x^��U�/��?�����ԏ;���e���	�_｟R"`l�F�U�7��]��=Y⁖�R�~7^��[.�e�B%6|=�t��/�*R26%t�.`"2W�ύ����L����X����_��e�t���ԍ}��bY�����6jE�J��2YV�@$
�»� �VW�$�����3��pb�����O=��aq=%�W&F�z7��%���j��4��1�;B�-�W��|J��]gC�EP��G����S�/,��-�-f�7��=�Y��ݯ�T�#y�A�]s�`к�裱�i3��\;`ͅ*�u����A�"S�E�&î�������.�Xqa+@(��B��)7��}cR}U���\9(}A_���u�+O @�P���'���u���Fx�jmq@c�m��#�M����&���|�pK�m2�/�T©EOY����=��n�N��,�Uu�Ý��n�8l�-
��'�^���ny��ԫhJh�dxF�T#	�/4[!�QJ���ƕV���r?�%��Zr�#�������r�z4��I��q^/(����{mB�}y.-muG��f
�J�����|v�ˉ�2���ε<�))��PF�Gm�&>�����h:�(���LV=��+�RB�B�bȁ��܏�X���=�^���C��2M��2?N�q���mМ����u<��p�&/��Y��qP����+���$�e�`Xy��PqW$J��u����+T/���k��k�9,��x�'�?4e�2m����-�*�L�Q}aX�m\*^�6(��3-��Es�(&t5��K.H�2��i�C<nmeh	�����>�/����D��5��"P�e��|n�M�_�O�)Y�H�Eհ���o�}ݑ;OHK@è�!�\��$����İ6���>�B�o�� ˄ܴܹ��XG�O����w����cT�fS����C���hvx�)����7�D�ۃ��L�������<z+��u���[�o�#c�C#�)ȅ�����@S�ۄ�����Ak^��%,P��.R��*;O��~�	��7��F��Cx���I���է����OY��l5��}={����)�i�E��-�Uo`����.�ɲ�=�-����/X]ي{�Z7��Ϛ��y����`�|<�'�
i<KLU��1�j/�G��ǩ�թ��d��	�b�&���� `�u�־�W�3�avVm���g+-����.��C>���k]�8�TF�g"%Q� ��)o���R�e|ü$�����W'�V��V(�6As~��)�
w�$pp1���j��mgH�o�1 ��$J9zb{��ʔ��< /�����;��邾���d�Rt������^���C���JMN
v���7�6���h	���|���E�t�Ջ�H�����3G8����l�@�R/`�4 M��l,zT��2�䓿���sV�Њ87�z����3�*Ի�51`ģ�7��������Mx�>M�Q/p�0�v��ݭ�#?�e=탋X������:�\)����(iط�ɥî�H�N�^=C���#%��Ȍ�Ĉ[�#���,�T�}��ߵݨ���R�-�]���T7�d,�'��x���e҈he�{"o�5���C�٫�֎oԽ�Q3M<�6��?�"�^�F��[-�@q!%�Ń�?7�
uoBj�W����z�U���q�UP��-�ɛ�;�j��K�1�z��KT��9����h���q��[���^
��:CcNRQ_P���ag�=oK~���k�'@�4�8�/Y�5�^��a�F��R:.z��HH&&��G���e
'1�[j���b�Hc`�:`)8I2�V��1G��_��e�i��S�s��ِ����E��T�t�^�ms^U����=N���"�$�I^�!�Eb�"�I��:�B/�Pt@i��q�u�a4$0�?��}�m���mt��,�yT�b6y�`�^�u�c9r���#��¤��O��,�
Gۊ�W��.�9��}L_�>b���W�C��{��u0��(�"�0�����܂%���Ϯ�J?�{_(Xg�>��������!��JN����Kt	���~�&_,�E���SZ�,]�͊J[�1�#s(	�;&8c8��6-�n��7� FG�ƚ7�rw�Avj郶?�����Q?ق���p���Y�]p�}���"H>��\��|���D�P�d��4QA�b[�ܩ���adq��0_� �	����νfs*A�HLJ�#���t�ZB5���L�#G��i``#b)w�̛�e+/�{��h�'�-1�,ź�N�IS�O��"w��#�0�431Y�!�����47��eL���eݢ��9zVjw s�C*��ˌ�a��G1r]��w��,�6e���^�¹ö/��#����-/�&��WG4��Cs+�TH��7!k���p*�ql3w���ڏ�!�A�㓈 T�� �w�~�ȭܦ��&��Z0�����f1d��� `瓬����_�Baո��p ����E�|��g��&�lv��|uk���iwL��6�a�@*���H�b��$��Y0��4�
H��[
sȸ�����f�*�(Do����S�ͬ�0/���1=��Y��L��C����l-i�������AU��T�W�S��Y@j���V��Oej.�x��L�ߤ�P����{.��Z6\W��o��K2ilm��F�"�ߏ���>���Ȑ��p�W��?Aj �.�V�v+�Ċ_�b�!�?It����(*f��Ji)�ǤrM��#x�n�[�JD��Vb�$V[�;�KR��a�Ɩ�CW�ND�I?$�j�G�}�V:� �L����7(jY�@��o��x=<�'V`�:�5���-�Ǳ�r�˃�O���pT��?R��$����5�з���qg�2�^�f�V0�ԤV��@���	IY&Pk�O�K�Uv�R�p=	��m�U[:����̓�
L��{%B*L0�F��T���UGȻyÿ�X���m|�cʲe3�7��S���V;:�N0�& �Ο~�/u�6����#�e����D ̵2��Vhq�&k���~;C,���3��;�Lj)O��H>���mů�3�RD�L0����5�G/y'��t���U9������������s����m%�{vO4o�MVg�Gp5���q����c�T[]��!�qw�t�XM������+<G`+1t޷�/��%����Vd�u���_�(D��P��o�^��>=�~�ZI�-e�s�L :[,1c�㰻��0(��D��x3��l*��ǚ�� ��L��X���.$����q\_�)d���j$do5�g;^j�����W������3�o���0Y&C�"W3_���h�ۍ-`�Ā�|�/�,�ɔ�-	:'������(�0[���Y�$��4��sQ(��2(�A�2��><<-�뽶�暑#q�T�~�0��ϻ��D�|��$�Ҷ8�/�x�I(�!E�Ɛ
 ��	a����q��_;�@�D�v_$y͐\�9����P�>~�*)�)�@V&4kW�gr�>���
��Ty}O5��_<��U��J��F���c8�Q�)^������$~٠�0̾ ���*��+K��Z�]���8/Q��sb��\�a;R*^�wMz�����%)Aa�X�\�iA��0�|w�S�m��_�G��.�B�=�a����t������c���m�s�i�N�XClf�-1��
ЏfgG�%[H�fb�#��O\ݧ�����񾞟�S�s���D�f���Or~o-%�wH�J�;�³x���P�?�,�K�5mz�����i�[-j�6oUG�/|��5n� D�U�pz7���`-��<���Ff12Xh�Yz@m_�Y��Q���;(�^OoI�'��^���Y7�@0��_A�ۃ��& 	��+m�dVvL��y^��0��Q�eG�3PE��a�y=^���R��WD<���U�ե�uiJ(�H�`�L����}齖�+�ɧH�!O4�Ђv�v���;�"���LpD�*�+�Yq}����9�)Q�c҃1��, �ߣ1��_�*�2'.�oy�:��ݶ]��t�ֽa��Y��&�I9[��+w#��I��)�e�\HhIʛ~��,`�\��sZ�2�zMD�\�M�T�*�Nx��ekH��Ӯ[����RL8B˓!giQ֫Xr;�ߍ1�3����mg}m)�P�L���ꖞ��0� �K�F���V����}�jO9|��%E��Jp�m�@�O�~C��<2X����O��<#�
�D�,�lkuH�B�\�����=�qz��W���^A�C�c��lI��G����Zv+x}2˞`DǙ{,���F �4;� �<0���U���=��Fq��*�-'=�H�@�1�7ͷ�V���'����Zm�M�RU0�J�B�	V`!���'�b"W
�j��F�����-���wc]P�;$�>0��+.+�>�^/Pݓ%�h��bu�9�^�>���E1���S�a���6��@у� @��J(�	=u������.�E������c�΀zO�[��*�b������^~*%e�7��E5�N�Z�o�-���,)"S֜cF3U_{����@����a��yK����b��{=���f���H ��x ���,��c��e�v�S��L�g'l��Q�����c�X�I��m���r�̰]�o'�12|56 �O@:���0�۬!ݩ�,u2q[�/R����69�D����ɘ�0,?��dl�)�.R����3�녃�d�Q�l��_��/�N��f�t{�{ ;$cs�NØ�ˬ�9�k�s�ѓ��ϯ���ѴitM�J7	��C��$ٰ0�N�_�#Д�;�\��Z���<�9'bW���E��$��p-14���y�o��3�xM*G��g�O<I:~#=i��bNXa� ܸ쇴�Ni)�L�م���"�ʤv�Vʼ�>c�_y}��e�>����է�>��F��p��9l�b,D�Fk~9��7���;�qGl�(dqm�Þ�"�T�m�N�D-�Z-����4ih�1@�u刽�f]�e��#��'I�����^�<�"V:Wޛ(r,�>��ض�T�O�L���Og� ���ί|�$5$?����̚'�hD�B|H����wN�۰=��l���ކeJ�*�q�鏮z8�$�aM�sԺN't!���4N�O�1鋠$�>Pi�Ð��ƅ�a��L�/��z$�6�_����#����D�yE3���$��_���	e����DBB���5<�\�ڂ(���i�u)!����!�^���-kȵ���}1�V�����w��I<�fI1�Qb��	��а]�oz�:Y64����2L��С��+U�q�ڳt�2Ƹg!����&�����G`K��(��"R�x�zF`�i��FȇW���
�'O�H�e��w�d�s�+v/Ȅ���e@�c�z�+�T��u^y�?�L)]��լl��F�&b�qC��-�Fwm�4��¥�ଘ�OW�ޤ�s�X��'������w���ƿ�1���=R�֏<�P�/=�)�H�±[ʼI�y(�ĝA��J��7�R|4.�3A���:N����v���|�S8�� 2q�ݒu]7�-��wIMC�V����.����������=D2'9�~��fñcc2������V��%@@s�P�|����:�n"�h��� �E��{������.sYы�tV��M�F�{��9<]��c�w�[]i�B��U��Qn��^O"������CKK�0)���������-���l�m��#V�* �uħ��g�W��[��CN��&3o�ݪ� ��I����ꌫ�:��$VD�U�V2�]���U��B-)���E������l�oB+�3
W�L�B�W��A��h4��X���=����E�k{�8<�G��� +$��RܘXp% ��A��TĴG�x�Ɍ���JΜ4��H3�O%��U��]�w#�]5�S�ƙ�W�S���_�i��+d��+��Ga�&�H$/3u�¼|,IDP]a,��kc�1�P $��cX��O�G������Ԧ�A��Ѭ^��у�K�.��=슨cM<�Sglr���A�Ec'K��[vP�j'�݂m�,cogI2cfd�ʉrϯ@�A��i*=/�n�.Y�T�b�Y|%lV")_�@�m�̘-.x�r7f ��.��$��h�`����v�9�S���Uȓ�^�ra0<54Y+>`�(U2#�!�ɓ���<�	�i��$[r���{�i*�c�-�cww�]OO���6�:�lv5+zd}o��4���zWş�o��ȉ�E����p�8)+�\n��u,C�շ�&�XU.xc/��vG37m=�[��m֪��>���gK3t9��Z����3�m�>Ҍ�x��yʸP�w��{�S��	s��A�s�!B�p�O�M�i3�����ky˟�9:Y�d�Ab���X�q��#�AS��H h:b�������Ki�fϖ�H��ڗٱ�K����a�\W���þQ|-N@�pL��ۍ�%Y�V�����Ә�g~�R?r��*v�5^0��@ܲ�N|<��ɵ��$@���3�qEӂ���>�P�K]	�~��(�¸#���COB�E=���)�� ��	��%�4��X�;sL����`d�$X3��,�������.�	An�����qZF2��]��f���Dq�hڑ��c�����15�+?�xs􂍺m�V��m"�<���*���S)��;�o��|�W��h�蛵ga�7���ex�(6H���)h����m�۞�g�\�����+��H�Ž��h�YN���	-�z<�):cߋlo��R�*Kk�/78^�cI��{�6�rW��*��{��lC�����%����FG�	��z��"�a��]P�^�ڑj��<�;�K�1�nBE"�,�9�k7��;c����x;����p)r[��*s�Ź�Q&���Jɗ��⛹sۙ=��q~�̙��Es� �Vg������.���F���g�W@� ]�@��G�K�8����=����E>�7�JN�:T�����B���'��7�q�kG�ߗ�[E�Q�����^Yo�ȹV�t�����fih����x�\��4�1�qd����KN>X��U�l�#Aou��!9+�5o��s'����F��~~���:�ھ��!P��`^j/��Z��%��E,9��D���Y���`n�{k��Y�!�J��>�P�����T�'�ݼ?{��#6���$[���� BҢƔ��I�B��n��}�E�G�@��y~��o��
%��a�D4��^�\ךέ*�E�W�j���x8��d��|�唸����t\�8�z�Q��M�Gj�.9\�:�k�Rr��̚.��j�94:ur@z�x^}�SlEMsJ�y�C���K񽴃١:ż^��"*c�������0qв�XT�x��!��.3SJ�E�N���~�{#���%޹S�槙��Z���iV�Z_<�'5Y8"E:�.�x҆��]Ju窅/ގ��$`'�&G�`đ��'C��9�@�tvmY0����ڡn#_�I�$�ť����}|� H	����t����!��݆_��F�f��sI_D�@�2�F9_:|�����X�*��R���#�C389M��sL�T���!xӆ6�S04܊ec�w@���N�k8U��K�{|ēP!6����ۼ[���7/'U�_� tk�	*Ri��VU��S�F��	��W����(��xUg�?h�K���jɁ�[�.T^��y�d�3S���~�飒0��'�I��w���i�|\���f�ϕbw�4Cq��#m�z�3D������ �V7�d���"߅���Rt�Nd�U���� 4K��r�V�F�rv�2͠E���m8T1�Yj���(��#`�u��k�%Nm�6BO����%�G�m�u�[�#_G��?a���ż��"0����%Y��rpc|lGx�/&6�&Nϗ��.iÎ��K�`����`����<ȏ�>��ݥ�k�z��f��{���*<§�HV&��vكB�a�5S�* 01.�2��O.m����5'�O�B���hm>n���-�aCbD4cS��ño�`BS��$pcxl��nG�=(ь���t�e����W��� �AY(�]-$W[8��B���;rD��bf���F�D�GԊ!�S�	M��[&?����gf�)U+��c�t\ez�a>�˔'JK�3��T&�&�&C�	��0c��x�	W�Gۭ�#&�M�&�S��x	�� k\g/l� YmA�) ����Z��rt�k��jY�F�Z�P�_Gu&�u������ɼ�we1�ݥN��Zn�y �j�@Pv�n��!�xB��ǌo�A�7l��{� V��� ��<-�:�x�K��r����3�^^H��� $�ނ�a٥Sc�c:-�����By �w&��Մ��>:��|\A�s���I_�C'�X���CZ؃?�����9��_D/
��h�,i�E�RM��䣻�\�2EBʌ�4�}�t��Ƨ�^��k�+�p\�*��o�%�����x�kͫ6/5�G�ud�c��[L��-S^o�t���y����kϫ�ΆƳ�h,���ؠWpis��y$O�LҔ������s�cʠ� �ȯ\�;���Q��R�G닰�(��`&�cD�-v�pp������q^gl�k�����!C��Ѩw��t�b��{�z[�z�1=#ά�4<]]w��d@M�P�e�U�9C��1����k���"/�mtr=z� Wm���/����ZH�w��|��[Skw��71����?j�,ck��}D}�K�)3�W���T�{'��lU8XVq�8/����QfU��	�x��@���_T���hnX³/
+{��)�������%>�r�-��zU��@8�Xw1~�HJ�1���縷0�e
�p�@�����R%�*D��
�9铯)��:�ȥ��)ޣ͎t��넹���<
Ξ�0D�����桟�VB��a5���[�{"k��j�aq+z��1���#��Y��������+�3(.H�
�t���èq�(���$�E���>�Gm�4���BO�]��F�&�mGOm�2���FI��f���`.Pːzz��<�M0䲅�a���;�׽�.�f�pc�:4��e|>v����<�����)�n�AT%.����ǰc\2�E@m�]=�2L�F��
��	C����/#dե��>����l�l��%�q�Ee�B�~���/U�;����D2x��kc&��H�&ƛ�8_�Ԁ詗��fCc)vw�-Iv���V����ㄯƖ�he�j�S�Xtre�=�̊�2h�]h���d�H��aNG�M}��Ug��	C2�0���ȟ\� Kn��{)e��Z�e�q�O���o�N$yn�hc� )�Gi�{J���<��!s����*���e)�?L����^���_M���#�v1�L���D�A���X3�:��p�J�@:_>{'�x`�@ܛ_,�֨��n����9�OC�sK��������X��A�f"6J��3�N?C�pUf�!=�n/w���!=	��1
�u�����o�#ng���N���yXGj�`�����qW���-r;u��3�t�q�.��7�+k=vހ0u��]fʃ*���nO56���yk~����eӃ�?���?�u�I�-��i	܄ȿ��s��jT\������ Ś��u��x��˒�����ݩ�򏣩>�8.�qϬ�f��ij��aXu*��WP�1�� Dh��%L76q֭�l�@�X �ɏ�K<+ܵ�4k��s��Ix#]6�Ap�`e�k�I�)qڪ�,.W*��{3C>´�0�$;���'n��{���[������H�x�f��/��~p�m\Z���_�`����e�{FG�wc HLl���x�,Mw� s�����U���T�ޥ��D���IyD��gq+[}QF���B�g[�א(Z��h}�B����7�,�QC�!�'�
x~�uSHd����u�qh+��Id� ʩ�H.k��룵&g~1�`Z�v�VNz�!tD�P
4�{^v�V�����Y��vA�'�2�<?3r�קUɮ��o�����_/�/�
����6g�-K��%�����'�Y4
0��O.!�k��q�K!�&p������S��Bm��ot�`D�pΉ�!2��3�0�%p�?�Ae��i/�����&�,a"Ao�)��z���I��Df̏����:-��e��Ş_eԕ��/ҘѮ����|\��M�G\� ��Ó�zzGHFV�U8��"�V�-���n� �����\!J�#���z���'M��KO��U�bRW:��߅G��su*6����EsN��P4� ��'o��	�i�譼W	(�Ȁ�wFW����W�}�uG_�������GҸ������%�֠�̆O�/Yo���n�����;YA������) �uё�o1����V���k�j�]���a�:%f�ou���m���(^��5C�bS��A%�qJ���Ӹ��t�d�+�.���%jAB���H�u#��֌�,E֔	2���we�r�|��� X� ٮF����$ZR ��
g>��t��%�j���ᮐ�1(~���<F���HN�6;u��CDn���{,l�h��qj]Yk�N>,�܏�%����s`�䤄���Y`d�W�SF��+���P�ň�`�~4���Um��r	J1�����xc�qq��[%{�^��<�����5����)��Fm9S���qxG��{[���� ޤo���?6V:��<R�l_d���cȁ��0K��
��9�d[+���fM�z>��9�ՙx	���7N��@Př0�rӬ�j%� 7�&W#z���;�EJ�	<}L��^*��<M�g����>���v����̖);�[�6bŗ�w��x5����)�sje"���s�/��kp�W��xzD��m!����R`n %)���>�?�q���D���E577T��A�[/��i�g(������q��ϒP��n!@�,ΠC�]J�J���� E;��}f�O�G:���l�m:Q��j4Ӯ*婯�Grq��V�)�EÛ�D��6�n�M9�q_^��yq-���UI�h#l��\�8: C	�5���s�O�����Ҧܛ]!��{}���1)�tO�a�����𔭌��y�?(t�lSB`��GI��
�xё��F�Pu�=�5R��S�K��y�A��>�Ch)��8∷r^�{5������!�6�<+K�?��W�CX]{���r�w�a��`�!膾N^�q�dW�,&ŇÈ�6:*��O���{�`C�e��A����T=pE��j���,� v��x��ݷ�������BB:Lj����N�wю�����r���!���)ؘ���"hd��Ί�k�n+�@>�~���B�T��CmmŜZ�^���@wX��)��E�@M*���˗}'���?��s"� Qh�ߘ����)�Z��+8��F�����}�\��7��4�k\�!D�V��)AYyn���jU�Y�f�Z��F�`8 M��
����Veo o�_�|��^�3���XQ�M�z-�&����p�ґS�>�|1S��et�����H�?��b�YH#�e_޳Q$2A���QX������������zr1?�օ��w��ؤ�J��U��z�Ĝ!J��9A�N��z��?R�ZDb~��Z4���^���ס�áɥwib�����]���NIM��lu°M�09SMﺤ�!o�I^�X%ƛĕz��g�	��Q>��;�M��<zQa�[d��,�*ۛHތ��;�v���s0�Ǉ�%$�\�r�������x�8&'v��5�������,�	�]��c�e�(:]��Pa�'����zhTn��6��h�Lzx]d+"�֖��)�.����,�U|�|-aǜ�����Y8*�L�l��l᫡" ��LM1բ������s�nu�<��ǁ�ӂ��T�}b�m�ա��u�r ��w]I�DZ3���-��
o�ry9���d��e3b���s�c�$��e������be^Z(�H��C&��fm,����&yۀ
�b�����[�&(��-O4�6C���XF���}�dP P�W����mK�4��kQ��4�b����ʥ��N}j�ZK�-�=���m��y�M�RR��]��L�f+m����"���I#����Tӏ�}E<e�(��+�f_��<0$M�72l�K�_'��̸��}����g�4����*������A�>���E�l@���o��dF�k�az�l@����x6�����.���6}9�tG��"x* -�t-��������H�֠�-�c� ؇��M���b�E�C�$��z�e�n�uտ,;����v�J�.
6�D��,9Ǯw�O��WD�_y�e�ho�|PVvC]/(BSB�+�_��i���^�&�����
�; nl�i���fx�>+Y���W���Sbry�)�̒φ��1zG���TF�H��O�L���u�8��jdy@:�i��2�\煿�	���_XB���&n�9@�gg����G,~Vtt��|��%�	�d|*�k�2rѯ�U����j�fq
�j�&�o�О�`�F��N;:W0U����e�����j��JDsk��c�Q���j>ô�ŝN\�dixWoڲ ��D�r�,��;�h��Qmr�oJR>%���M�18��w����w=����_�履�Ca'@^!��n�B�X��[��?�KH��Lh||er�a�Tv_�Dk<�/�G�τ��ؕ��Ԉ��tR^��5�-Ŗ��Ey���kȬ�x�g@�����[Ag�2�o=����!�Rה�<4|�"Zb�F:q��4<{��XTs����K��Ћ�.*�}�(Fk`51�����bj�X��H�d�ӫWY�QfB���7 �߹�n_��Tz7̊5�՟�؋9��gg�S�H�dH.�-����+Cb1��ҧ�q�6{�&��I=1><\gA�q��uْ<_���{�bQ��5���ߜ� :/q��βAo�iX��6L(��`U���rU����-h��e��g#u���^ol���M�C����2�I��eM/�BߢUIIJK��q٫k�l���*e�їI�m��Bѹ��
I[⻆�6o��LY�{��,Q��Թ�����d_6����͏�5�X,�޿E	�^e{�1u�vmI��ư�����]�"�#���T��ǲ��^�3��Q�v�gۢ��z8��s��X�W5I�IYM���nA��2�˄Y	T5u^�(��$vl6�W�[j`���P��|@�����wr�=����1�]�Q�6��p%�f�2b�*0�n}U�n�n5����$�v~~Z�Y(Gl�eL��a�s8|��=��|�]�.Z|�a�����S���m�4?���Q�u*�u	-� � ����3	��ٰS��?.�K		���[p����AX�JL?����Hm��e�ŀ'��M��2���$�Ο��zV#�.�l�?ג�ZR�ʈ[;��V�:]�lb�j��B�)R!���������WW��[ڱ+X�1�p2�4k�1�$�4�[`Ύ��0��G�c)g�(ʳ�O��z��z��\gxa��"P�M�y8�?r�o�Dr�,ҹ�
�ژs3��J�S��ej=�Uw!<#���"�\S\�}V�z¤�)�A&~��o)=&���\�l��.�a��7t�Ƹډ�V��5c8�x�j�����x�Tf�W���/�aֳI���13�5v7W[���>.�,i����*сPE&�VReC{Ro�b���P�Nޟ���bfM�$F��s��]���� X��d%7.v��d��@��0���4�u���
p�{b4�d�ݲh-�iǰqٔ��[�7�xu�Yv��K�V+�JE+�f��r��j[)��i4ԇ?4����pi�&yϭ]X-G��cdo�'�W����ƺ7U�޽~k�c��=���)l�U�1��x`l]׼e��Gs�a��0�.�߆��*p~�H���+�*���$*1�����2}��}E��@M6�'�����F�8�n���~�������J��΍B~m�S0R�!<��A�};���l�e�pC�Q����S
�4=a�:��Xڙ�����7��0��-cXK���9ͷ��J[��(xߓ%�-e���}�v�\�:�?p��x ?��A��Ǆ��I��Pc�Ɲ�)zVI6�L�m#����Úe9��v>�YH�õ-	=�3�0�Y��A���L[lU��է	��r�U��w�#q��{92�=r���K�|a弻���������D�+TqpX��M��&k�v�]V��N����ms���d-�=��1�q�rc?��W�5�+�E9J_�"IC."RýՓ�j���EPw��*6�Lՙy�e?�z�h�"�҈�g.�Co)�,�cR1���?���D� L�"υO�/�6�q=X���A�e_y�7��R���\mGu:$9+�:32b7M�DG�,b;��/���˅xP�c*'��m��O�t{*�rG6�'I>���
�~1\����ߕp�� B5S�UG���J��,����I
���0 B ��H����+,��Sk������|V&�,����Qc�CfoG���p�y�{XzD|��kԤvH
o��(��%!��L>T�_���Gp��:�[A[&�Y��{�_	.�~-�<�4��u�.�I8Q�O��B��k�q	J�s�#�\�n�Y+U�l��U��|?VJ%�rZP�]}x�R��]�F4�����/����P���͢uR�Na �%���V3�΄$~��H|�zK�U&E.F�/t�G�S{m�<<�K�Ĳ��Fҁ����^�#&Xht-,��]j�o��}KF��G�lkh`D������ܘ�i,���؄�[2l{���O���G"��:�l?�H�����;]^��Xl�Hݹ5︞ܢ*�_��W6�G#��i��Hm�0�� ��(H�<��0��7�xd�'�F5B�#�
��>9���Zy=���c8V�uQL�(�Ӯ�!�|�It���������O���irV���yp����T7��eW��J�ڻ�Dz3x�"m������Xm0��'������.9+rAZ~��/V%�����	��p�=%@�Y�� /�;d�T��р!��r�Lg�a�3�h��9�.���D���A���)�J�I�(Wi��xϊ�����fػV���J�Ji�w� j��x��P�C��>S��t>۽�c����?A���;�@C�����V�>�S�1܋A`"*�R]7�����D��@[�"��j�k�IJEC��}��l����^�B�(2� �t����"Q������0��-��V�z���?�����Ja^7��*o,�Pw@�5�5Ɏa6��BPW���SP	/�KR3kN9�T{Z��t�:�q��N�F!�U|�!5?�����9�dC?�~q��/��	Cb%�e#�8���7Ň�]� �Zq�s�W�R(�:��-7��f}���G�4����%�	N$r��O���7��gIE���^�H@+��et��w��kWW��I���&���n~y��Խ_2�q��1=�(b/�C����>��=\@�=Uj�w�^��<_��*�����Q�`d'���y��!W�6�g���4B~�6*YѺ.1�x���jH�%�6��6��
r9sN"��ig��$���S�)�2�E4�&m�e\!�-��sk}�g�d��U�cm�QPHb���ޕ��Ӄ�{o��Y��ߓC�@Y�U������l���q/9�L0[���{��딩��Ƭ�r���?�7c��*��{dF�x������&�C�����7\Q��E��<�`�� ��c-�w"js�u���T��V2�j��R�0�>�of���H�y����D�l�gN<�Ԥ�ʹ�����Gz*�>..ϣ�m ��c1�s&TI�M
]d<�1�t2yO�˥�	玨���}�H X��F�m��̍��+ <8�Ņ<�?��p�4b�f���!���I���Vz���3��d����uVE�O���&>�7�8�����h6�Jw1|�S����@��(���b�h��A�j=l��qͨE&�p��d5I�aÍ|H��v�,Z���o���@��i�gع&�P�p��-2�p�>�[��&+�x��M��C��#F���qK�+7ywkՂ�� �i����]G��ɺ"7s�t�ٙ��p�����
��/�1R*�v�������J�����F�*$u�L�{���|s���k�*[�]���":ꭳ�v��|��xl�੯���Hj��O^nT%�z�!�e��H6�S;������i�䅘�X;�E	-@k��,qnʈ��i�@"ӌ3��kL�w�DX�r#���4n�������I�fWf����}b�ٷ�g�LԲѵ�d�`g>���aqRn��PP���4tQ����s���֎���qǱ�P{/Qg~3�����ҁȑ�b]X��	�rŜzo�u�#4ݎ!Ǯ&t��Xo���!��}O"=ƅKBv�f(��o*������"�'�eh���c��d��R�m��gK�GS�+%p���[i/�:��X�>��X��Ω����E�����H�Kc��n4� m#>����;��T�G��rF���3�ׇ�v��c��\E9�D����9mx�ޕ���q�ޑ����Y��3�	�􊕚L&��z׫��l��V&�
;_�
�<X�M�Ҹ�k9�k�W�	Al�Q��mX���z����v��<G���F��b.7	gr�ߐ�G�m���Aq��+@����V[2�C`��Ƥ"���׌T,[���e��)�RH'�!�"�]n�D�+��bv���!�p��Ǟ��*/�9Jz2:׸	 ��5n�K͂�k���tK|W_f��ʸ�������VR���#�
B���C�۝�H<�,R/���a�,\�ox�9a���Ð�Ǯ<2o �>Ybt�\����bgd��F.ˇ��ZX���b*hp���Z�ֹc���V�w�3���.��I��z�����9/����J|�)3*#��2ޮ�F+2"��X�����S�M�A������[�e�e6���d0����H�gu[M|p�?�5�u�;#��]3W�c�[�w����	cn���=��[��|xŮ��5�}^t0�f�2�G������O=�b�M@��%�����{�W}V�P�Z�FsA�v����o;_C���-Ž�}��$����P@C}�c�k�@7�k���Ԉb��[�'Q}n%(�G�ͭ�+u�w��	��}&��<g+M�l������r��aޣ��M��)����~� �z�L���} ��(`�zF8�l��3!a��g�H(��~�^$pHLT��$��x���H��DD�ђ�����"*r�o���!n J|�O0�G{T� %����sx�kbT������&�g��� ��b?�k	���*��s��� ��LU���mS��_�"���~�����Y�� .�A�X`s��ȝ��������H��%���$J�&�W7`�^&mW��w�$J��z/��0�������]\�Y+�]�|��Rί�u��
��oY�U��瓅��U�I`gSp�w��7xyW�a�#��]k7�/"G�r�KϤG>s�#��َ@>Ó�L�����f�H�zi�>u��&���4�� ��K��������=�g�!�d�I�.v���;YAD�u�66�ڠ!��t$#�H�W������Ω�n��dn�,(��v4Yƙݲ�Zѹ�ш�� :�͊���`�EN�6�T�/	�}��|T��ȍ�K<��c�������%�*�4�k��'������H�"�C#�6�JU����Y���̏�L]:����E�"�W���$Q{��w۪�}	��y�~hJ�O80�0�W�F;������<!���R���(�S��~��Ϙ��P���2�G�1�q�C㬖UT���$_$�[q�o��;ۖ�����[Q�R���w��ax�����&�U��&=�����֟�S@�[�_n[��W���B(��l�j�*��R،�ѭ�p
�s�ZߥZ���}^�d�/X%S��l@�`l�uf�	*x88���f��Г��"m�5l�Zé�,Hj��PJVIz�D�Ij�ؚ�$�?�?�=�T3'�h�gj"?��;Y�B?���M��Ar�,�U@��9ٔy?8L�Ӳ���������vBL������T,z&�>_$����{���>Ζ{ǝ�V���'�1�u�Nh0��*�P��?��/}fVWa���!'I!`? !�߫�U/�:@ԥ~��q�N4�4R�L�l�� X֪ු��e��b�fzw�r>C�����
[�G@��ؑ�gC��Ч�'�b֭�"������DT�̎\aq��a�O!9(�^��8:�&1��w��s��w���a�g����^�늈"2q�&R�*y��,8���N�}=�fQ.���U>�WWa7q�H���(4�%`�LB��E��TՄ���o����:�dN����Ѿ*A+"�6�Y�]b~��w{F�������V����$d淕�&�朡��֔o�>Q�$�od �gHW~�gقG�I&h�D�Qa�܌��;ݤ���H�s=,7�$��������n@�8A�)���#<p>t�UU:��%2��w6�횩*�`I�q4�0s�b�����P�v�K�T֤P
�t%i�g��I�o5�Q]O�����R'(	��G���,�;��)��DT�/�Vץ�,1��
NY}�A� YԻ����T[��u�9�db��)f���_��7�t*�ãuШ�O�`���T�@:vcw`I��I\�@��a�9��n{[�(���3ݻ�ͦ����y��E��TFxWc�ZU=�ˎ4�V<c�y���k2Nc(�r��"�Q�$�Z��w��}!���7�:'�%�{����I��z���<���T���z7��&��M�
�@�(��M�V)�!�\/R�t�Ck�?��4����YE\:�&���%��`"p���qኩe��.�/��I�y��E#.������d�3.����Tf�t��Qē#��X����+*���]\�LǦ�>wk�J��Κ�+�P�׊�~Eg��J��2�g!�)X�wP��9S���(���Z^���Y�����	2�	�!B��+��\˯\�o=$�s�yq��&��)<j�
1B�IۇJ/M@��u��J�p����1��@�W>_b=�2L:�g�#�>�k]%K�*G��h�~��D������Y{��]��؉�.dg��*!��&
F��:[@_�4�?�E^L��1PT[k�B�����R�>^n#T�<D�2�w������6M{*	� �pv]B�%��Z��6?������׍��L�p�P��;���hgKM�2m\��2<r��~���yYy�6m� a���Mwi^>g#�=����K���3�T����R ��n�Z���h���]�+s��ΟF��܋�����D��2n>IP�y&xp���]���-�����A�p~؟��W��J�����
`��ϡ�����f�+�{�!��ݝ\ )Y�K\�~'$���)ETgV��}t�Ekn����Φ�<v�Ϻ��%x5T�tW'� 2��c���eFv�5�pZ��ӦU��6�W��%�N��<_��� �(���J�-�sZ������߮�r��#%[B�q�U;鄋��=B����_u�.�[̘��O��':�U�t�Ɠ�.N�͎B�6�3L.�y7��z�D�;�#�:	%c���@J@쳆�GS��ƌy�d[\�y�KXg9~����'a>*,�p\���?�﫹�Ԟ9`���N�-�&5%�8��)�1O${XX��rc��4/�H�r��,lA����`UrƻRW����~R��zy&ƽ��"�:�����'�6����]����M�۽:\�r��0ql�X�^�; �Oy�q��3!r����0�<���nЉ�8Z�C�����E6VX;Y���� ����t��;|�o؂�<#��-��$�e7�	���DU�3����7�O�{(�&D������r �eQ=3T�w�`���_G�횑v�=*��0l��taY(�)^`�
.��P�	.'�G3���%G1�K�Ek����Y�B�k|!�C����i���p0�+��	|#y�m��!��F�\��NТ��3֖�CZx���nN�a�1_);!:��4�#�&m�v��vzO1�s�m:���$B8S(���®�e�L�4�)+^h,F�r51��a>	��L�K�d*�������/��#��:g���yH���1��U���U%��1�����	��f�/l����/w-g4"�X�r�k۾��L:�B��9ث��"�ws���lx{�s�Bz�J�j��A��z�^��J�"�.7js��߰s�\���)/�� 2��K0�B?�5~�&�k�*����q9h��,��Z�k-e N-���:qBЁZ��K�j�9DJ���D҃���O����)�D�����Tl\s\�nc�]oH �a��{:��.�
����Z�������C�'yw�bx�wu��v]��X��'*O:���O}z@��i��f�g���C�R���uè��>�ň�%x���&Ԍ��!�U�&ѺAޔ6�;�Q��E ����dv�7N�F�|�vI)���c�΅�d��|T���"^�L�B�9��Em�98"��;��,3h&4jY���j�|��~���a�2PB�@���fz�� �oC8�@�c��!�YY�U
��DFk	����//��_Ѽ?S�}~�����Ln�T)^bjV��/�^զ�C'��Gf�Q����`H`7y+��,�����!��#6oBc�S12c����0"e#�o��[�s_������@��7wr'�Pʓ�8o�ӏ]�s�L�=C��9A�_D����ܟ���u}�$ݒ<�c����8Z39 �2^���Jf ?c���e[���Z���֗�-?�O���u��f���:����Lx0�&<K�aڐN���J:�Q.l����##�\M�ڙ��1}k6�Ys�i7:%O&�l�N���&�e�o	@��7�f���<�&��\�r0��/���4Z�089sV��'����&�ԋ�D�8�R(h�R�G(<`�bEZ��ni�iE�F��<��]�������u����Q���PG̣�轊.�:��a���� 
�=w~��;��Y,��5%@WG�1`���0�Ĩ���ef������M�+�Lg<���S���<I�:R��'o�|��'����*,�s�b�\�ɷ����1��
��i��k�M#\�;q5t��߱0CR��t��j�W��$�la(|�,@�M���Ь��<`��Jީ�@zNNS�KP����H�7�a��n _h��Jp�92;��]J�ຒ6��U����������u�@tT����O%��i��K�x�В�R��ߐ��A	@z�������=�]ݙ1c�E<��y�׍�'�Nc,e={�w��-����"�8/��̶�\�Ձ�3����-9o�ʜ�'��LȭJ�`C'_�s	2'�+�s��r@:�0��b���]�t0bw>�qA?��B��� �������ӵ�:����{�����\�� S�?���%��B�G���V��m���X����@��+��Np��ܰn�^(5�F�l�8h��='���U�;rڹ�5�HѵŠH%�.=?�m*��x`�M��>o��y�;��8�g�z��Ȝ.<N�7ƒ��DtSPK>�� 2��Ì+��$5��i*/�C;�ekz�4
�Ij��Oh��-��"�h^mU}�/o���j���O�t�O����3��ض�ӂ.�\���fѐ������O?�i͈B����	���~-P�ft�v2p����З�����s��d~S���f�s&�R-X���
f_J�/	�a��G�D0���� eP�� t}'4��6n]����Ծ7~6�v �N��5�IlI�y[S��J�2Jxj��L�o��o[y�ٚ�T-�Q��u6����.��=��Z#�R�dm9K߉���RO���NvĀ+�z8�ms�z��E�����
��݀�\,��D�K|9Z����W�I�~1v2Jˏ�B�X	d�!�<D�Q��M�x�gJ��!{*pႤ���C`Ć�~{J��&�"��O����w0f���n2���a������iBI+�����t�R�;���*�\����9�j(�綔��@�I}�C;!�R�z'Qmyȅ�H������0�8����8_ �^[�gY��3����N�%w�3��jov1[r9G����%���W� L̉�M-���x'ÎIJ��u�i�N��sz�݀�*�
FӲz����S��{g�T�7�M�ҙT�U�~�=���!��,�¢PE��0���[5�I�IO�!��^O���s���9��Ma+�3�ҝ���:�ny�.>�������)<�wk}f����|��{���F�R�dsC����!"Y��H����I�B�?�ŲGf���z/�h�>��.x�np����WzT���~bU�[���7d2=�l9N��.�g�����|�~�Z�קϫ�`�U����K�	��^-�h}MOj�u�}$��M���fٰ뫭�a-ꕔ�u���G�u4�R�Q�:��_��*/�x��_OS`���ލH��(�4}Ϗ�vF�"��t�9Y7���uA�ؤd�FP�K�
�,y۵ ������y�;ͺ��i�(����..�CW |\��-�nG�l�6g��?�{3��hf������!��́SQe�
O��74 Wg C�>}3���t��6ʕ�H��>i�����v�#Y�9r�����~���U��}��H�S9H�ԡג�����F�إ|��H r�|�L� GuV\�|Q�S�����b]���^��D]�M84�̽{鿇���a������EWR��\|�O'鬹C���,��u1��R��9p�����	��+��O3��Z���S�p�1QЇ��M
����W.�5mєI�2
Y=e/Ѳդw�u�%����3�ְ��ecb�*�@D������Z<����� ��� *�^Ng�[%��i���5��^�*y���N\F�I�G �ʣ�3�g���Nn��F��Cbf�W���& �>��/�����4C�=;��d��حUo�!?B� �����e-O�(]��I�N�Ӑ>�H�(E�P�Bf��|;u��I�����?�@�e��GRĕ��VP�%_����>һI��sB���jM��R��Pȣ����w�1M�U<Ҫ��$UN�-���Y�+akfA�5Z�3����w�\S�g�h��"�;��"�NH�����|v������v->Q$�Fd��G*��ie�Jd�-E�є�q@E:�ܕ�s�c���zO��9�&m�nO����XG�:3,�qc����"~6?�����G�A����~�۷�n)��۹;��<>,YPk���B�L��n�ҿ;��A�T~Ah?g�UC Y}I�M"k̚�t���.rz�Ь4��#�靠M_�/5�F��y��ݨ�M� �Q���D4�W>��L�a>�HA�is,�o ��8y�$�I�P_��h~4�A�&��

Ԡ� LT��1�ls���-[f�ڹwmAZѭ�<۱�p�MA`�����.���M:� ㅉ�~� �:N&�l��l�����jN>���⒤/��3�/�Q>�]��z
���h3�T�A�G[ʖ����@DV�,<��-g� ��I�%Ue��&Q0B�w� ~-l�"e�'����0M!��.��;���[9k;��Vݲql9�����Q|l���j���.�4WR���Ӌ�v�g`��.�^�ɧ�.d�����E��o��[�PE�C��]_���L�\�(��΢ȏ�$\n�U)Τ�ԓ�*��A��c��X�j���?=ô��|p�Ԁ�hN�dđC����CF*��}k�Nuau�M;#�!Kp�������#�1�-�+�γ�;O�&�z�j�p��oG���@�@kc]��W�Z~{?���׼�&g�ù�g�]M��#Y��=�&4F��6�5��5��J(��.t��|"RTӜ���F��o������ҕ~�E�z-�w[�Ռ��{��۟J��,X!W�-��h��w��W�C=�0�?�F�DZ�M�CC5��ts^���i�0ݞV0��}!��[���^33�b5ی,�v��]���Mk��鸰K��Z�\C��<��~��L��%�Y��(�Z����\��[~��#�͐�f�no�9;�F�*�0��]�����h"����`D���s�Ԝ�UlFh	Y�x�m�8���"�� �a����Wt��ĺ�kp�D����PEw���D���p��i/��;��_K��4��FS���Yz��3�#@���ȷ��9he'�91_����/����f�CkM��^|޳��{�ӏ�87M�굑��&Vb��"��ߵ��ZJ���������3w��#W��K.p���K�R�E�#�>���Q���I�����&�K{@;O�P���`
<�����{@��$���yEܹ�����'4�Db��Y���k�$+���1�S���`"9��fq]�XD��M�|VB��}1��_���9,���O��d7��	*!��zO�
{�j�_�8��JF��r�m�S��#�G�[��� :j��x�u=����;�^u[G�u�
1z$at����vTX|���GQ�>v�Q�%g{�O�"|��k��(��YO�lm�خG��x"�S_��b��U@�쫬w<F*4FHM�{�{y��m�Dޞ;�s�6�ͥ>8�*�3	��m��^�I3�߽���� ��#I""RC��RE,m�����_:��Ք%E��Ud�kK[����+Y��jiX�R�f9��oʚI��ᖺ鳼�PVN#��.��4�+^��ӟ������ɼ�7,@��Szբ���9_�~L)�.2�����f�n�P�#[Zg��SanXr��.���t=i��?O#�9q*��M��B�U�0[����Yl:�jzYI��a���}_��$y�K�>mf&|;>.ԥN6�m�`�]w�5ϗ�.���	�0dڣL�����BЃ��@�6.��7l'k`�������t�
E⣽r[�5LykQͻ�+M��.V��V \M�sC�Z�����z�FI�RI�)�q"��:��H�_V�>�� ;mH���o��bv�Xk��Bcᓾ��ǣ�k�1��|�ŻaG�z�r���x�SJ�=��$�۷D�S7>�]M���3:�ق� Ba�v�Y��{����<P�{��L��GՑ�,�B	�����5��	��ހ��PQ�:k�nlE��Rx7��3�������1������h�������\E��mϋI <Gn��c60�w0<=0�2�1S��N-0l�d�Bȩ��̴W�6t��[I� �����J�ä�S��`j ���4?L�K���%��~�/��J'>яu�	�WVp�Q��Ҭ���.���p5�uJ�*�>[�N~��}d�ۑ;U�M_�LB��������z���	�u9�ڡV�8b�	�H)`�h��5/vmV��dA]�6�;�q��F�������TD=r]�F]o���	�
�/)�V�)h�x���F���z�8m,�<������_b&򇤁9xh�� �_l��*�t��t^�Ճ�����9��8���ս��Hȗ|��}�4�U<u�*Q�8>�iW�J���s�(>����T�
�9 �p)(U����������	Gڑw�"�.����,F!7f����+c�;K'8xf$��QSfbތ(E|��Vj6P���lb}	�O��c'��j���"���B �_#��'���7b��ڕ�O0�0뢽\�5蟸�%�o+��E�4`_!d����'�ZgK:~M��I�g��\m�°��q��;�NTG�F�7�΅=%2R�?~ ��f\�ŘZ�q{�w�5R�	���dQmN���?�<-%uk���ޮ��dAN�g��ð$�}~�I�sl�7[�fU�����T],30���c�6 �0Wi��3�Y\�A�z9�J�]�2�����!�6�T/~���?�	�WF}u�㔷�ذ1d:I�Z"����D4ۧ����썈�SB7_,D>;K��%&H��e���h���YD%�E�����M�?,�K%̓���[y�<+ؗTGΥ��U�4ʜ�Y�}r���� ���z�}��q^һ���L\�A��oaz])&=`��k�E��+�~x���f�~>��>#LD��/�T+�Ӂ3�O��@تS�n�RNZ�u��/ÔX�V�}��S����tlZk-"p :-֌f$��Ȭ�O������L��$a�y��	��0Tl�K2EQes��EE��b=^u�p�N4�(%�z�u¡���2ֿXw��d�����\��Og	T��<����x�h|V>sT��p� �3_ݲ �G�Q�����f���1�i,�dY'�hWr6V%��jf*�� >��/9��r��h"���#��Ǻp�OC�0�-
���·��U�\e�(�]�BS;���#S���"���&p�Lo	 �����43�A??R�\��Ɵ�u�+�%��ح+��y�ˢV�yu��}��Za��^�m�#I|@�k�>ӛC�}�1>�B�jZ���0�8p�_�^�w-1`(J|.����m"v�-�Ȉrc���ʠ)3sH�~D�J�$ጃ�t+�%�\r�������5�v������)i,ɏ�9�5��"��,������U����D0	�r!�	��0.�]>i�ݯ��K��	���ώ�І��H@�x:H���Di�R��q�ֆ��SI{E�a����o���h&�t�|��ܬR�$5V�~i�T��)J�	@������Xr�Q	�\#�*�#�����ݑ�6i�9�`��n#�:s���Z��<��klL.po]�#�$B켲��-$���:<�v=����QA��o���oh�	azjr���{P:��<Qy@E3�d�4�S���`>>��^�h��$\1z~zy��/���Wz��h��ROP5�.#4YYƧ�^�Dˍ�[���m/]{E���q�_tV�`���p+�~MjE���,��jy]�$��뢫*·�d���q:�r�V��A�Y�|`'_����4mg��%�(5`�[��@/��@R �眣Ő��Ug"�q�C��Z5`<�w�u:$T��ۅf�Z�<*V��*<YAy�����>#g��|��i�6��%^V�~M%�z2�_�����r;S3���')a��?��nٟ��([e�g]��t0V�)���[�'�Xz~�����4�7�u3h�<���7��_U����NNan�����Ǡ�^�l�&`�WX�n^Ã�W�hq�+�BH��a'�~b���*���k����xz/]���s|L��=�h�//f<銌��f��x�>����KG����́=M%��s�I�LNN����t����X�H�kեcț���X;S���Z~������ѩki<Z���Ad����׆���du1hJK�}���58��;.�@��љ��<:��Q���zXޏ�i��w*�D �?�3�|�G�G=`�̪s+p>X�-��V�Z���?n1�N�7�kd����&�AY��*¾y���#���#_�[s{*��@ט"���2��7j�a�cr��7����j�wCs��SZ��)�������ݗB�Sj�&�uze�S.�җ��kq�=�=�>}�O5�c-�g��10(��s�YYh��A#r�%,�l�)���<j��C�MbxVtK�K`�h��T����T-�ܣ��QX��!�E� �M%f��U��t��~�'fK��N�R�����aM�q���y�Y>0}H���c3X�$bJ�*FEW�8s���Vҷ�.^�;��gĽ�������? nMta8\~V�t����54��5���V������U��\Ѧ�4u��:�Z������ۇ*�НJ���$�-��M�̧Õ��E����	!$�ʁ@�X� ���	?��m K�En�d��s}V�d*ED�We�Gs(�=��Ҥ��wy ��k@������l�1@hn{<�P­ �.�@ti6Y�;�����N3�Z��_�+.@#}7_�O��6No���Te��bG%@٘'��F�-](_.��;�p;��{*��h�윛�Ě��6�Q���ON�=�xC�����<����,l#�je4�M�Ӷ�@���.G���Ju��3r܋0�Y-�#_�	&���?�m��D��O��N��W/��G�@,�ᕳX;���B�L^��m�p�
�H��3~X<
���#��ޣ��`�f�[/iX܅<a���Hw�\p�s$�D��`��
����bҖ�"ڵ�ɣ��Wd��	�W��iO�w��@�́C,�>U�i~� �3�Ha(��-G�Ō~�6�|V�Y���p�Y"~3�FO0���n�s����4���g���u����g���z=��07`��c3�������
'2eh�|j8h�qF�ذ,�2ۡc�=<'RF	r�Y�:�nW����B�-qsut���Ʒ�4�r
����Az��B�Q	�5:�|L6�w�t?ڙ��|�j1#�n��c��w�v(:�v����:� �8��vg~HRI��E��Ag����5�au�w�,:GĜ�����'�0�SFJ_2�ǥD��q�,yi��٦-:5��|1>ް�,�N��8h��x���d�?|;$k@�T,�D���
��1�D�<I(<���Z�Й��V��[�8��|O��G�\		�j<��j���ћk�� f��MglR�׌T� �*��Xp�pq������z��K��gj���lt�����X\���h�~���98�
��B���p���*<�N��eu�T4.j��&��R_�����:?F��M�7uAA eSA�7|O-�am�/��-P�b0�tӂD�
�_�_Dm�Cri�#�)�Y���j!^���K��BuR�K�_H�{	aA�2�]�_��05��z�P孴��t�Mw��'���|�
B��M��E�\�v����Vz�ȣ��>��4��7S�jh�)�[DTa�h\��ɔ\�m��y�^v�G$��1DJj@����,� ~�]a�!>ڼ�ɦ��_��"��E��o�OcP���>C��$���bDd{�w�g���e�أ g{Ԗ,%;�{��3N��״�R��J^����n.~�8���̴A4,̑�j�'b��??�p�f�E,�Q9�y�Q��J�t,���́����4]�(g&n�'� X��i��y�H�|���2E�Ocsa��C'E��4�v\�z�l9���stitOH]�����������L�1�d/M� bP�K���;����L���= ����
��b�2�M�n��^��b^F
ƈ,����~���	�T�\��{�`>z��d�W�l�5U�!�&�� �4��T�6�lwN���z��OH�����hW�_$ �����p����~��n�TR�TI>��N�H'�u?��B�����v8���~5΁���	�<��G[!���{��]�[��-�x��R?�_�JoR/Zhv]�8 #�"��u�+t'���
�'��^�_(��遀�ϖj���������r@�a��Բ�*|��'�|��Xr+t�G��j����JŌU�#�[љu�FI@:5g��bh������bQ��a`}�0�`����f�F2y�C�u8�f�)���\���VN�(�j�A�"��0�g2 B,R�
 �ȸ��d��XD�P7��&��``.�T�er]��b0��Yѕ����#8����x0#����qD���+�խF��{FׄB��!N/[.p]ns��V�Ȃ��LP,+l���$ts�����j���
���f��>}/��]�ԅ����L��{BxJ�yr���wٷhW�dJ^��W�e9�W�	�H$����dtt6.!�0<)&J	[f	fe��8�N�M+������X���43on���z/L�4�+O�է���ۗQBK�y�L#�5�X��Z�nhg�Ebfp��O��=6�p�*kֹ0�Ÿ�!�I���|C�����.W
�����ǻ&�ـ�_�K���yI�p�˷�	���P	�^8�c}�ǓᲟ�j��1mEc���=�b��z��B�*z�?�����O�F��&F�(��C��B�H�z��go�����6��J���qA��*	�\qe�͂�2����35����x��·lF,�._�	����� ��(�vG��ş��m# w�9��1�e���v%B5T%E)Cx���%�t������0G���%�8E����zTh�GRI�2���y�� *K� 0���,�,Ia���4�Q0���r���L�Y�q��6��`�b���n���1�������PS)l��udO~%�n8��(ģG����0�T&�%�r�����e����8]�t������d�� lk'�ޚ�&�P��R��Db͆��(ߑx���IY2l6t�����MHhQIE+',`��kB8��ݵ���Ȩg��|�2h,��㢇�h]����}	�·PČ[{��>���z@W������� ��l��\(��'{ڗ�����=U�JڕjRX��ѓ������x���8��sm(�-���v����=0�L�Rn%8��ëO��Hh�v��gγ�k0���\����W'=�jb(\�?l�W���ݴi�傴����^�w9~�r<|��f_��\��%����+��Z_���^��/k=�O����a�*�7|u�C�<�D�Gr��}��C3�@^f2!������w��c��Ȱ�U JW=Ѧ��&�p`LO���'#�Yj���o�mz���R���_���*�٧���$��\&<�"�u��+����a=C������'Ja�KƠi�$�B@F�x�&9M%`�Q���0�_�xG�?t�[��*7��>�||>[u/A���xC�f�H4�}�FOi���i|��RӬ=�	���j�P�����\3��'��	,m��a? �)]�n��2�"��!� ��:�|�n3���<�)a�b.��8H�u�,Y����Rj  �&⠼��K���W��|�2:�4��Q�J%��������E�6L�>í�[.���-@@q�Ͷ�a��|�p9(�=ڜ,�E�:rF��$�3[�`&���9�e�� &ӄ���
�O��N�#��h���D����P6��M��Vη08TQ���O�2��(,��c�#��\���>�Y�Q|-��e���V�0\��N2���������5O)�ڲү�_�SRE�,5�)EL~Dn�.O����.Y�v)7k$��!�?^zD�5��n!?gZ����J#_8h!�XEj���+[$�_/9As_�0Q��u��������_}�<��u�tQ��l�Z	�]s�"�2u���5kv�	�ʿt�,�p|���Y�I�=� ��d@k6. ��❬92V��ը��M[����a ��d^�#�8�"�j�Ã�L�I��Ɩ��"�^3�Tҷ�h{�C&��r��t�&d�$�B��+�����{���B�ٱ�)�ҍ3o"���������������]j�� c�υV� kO���ݘH����u��i���R4��%�}H�Q��}b����"�j�į�*��u9�KT�?���� ���le����+b<��� q����z�V�<ⷠ�B�u�����'��H�ĈԄ�Ji��づ�0dB�ԯx� s�W�]6�I�'(ȍ�0S_Qk/r�'��vA	9���*4�E�!%6N�kU{�ʲ��q@ÜҚM�i������:�Ú��]Eu��~w����Fw�U
;M�	5I�����zk�l��&LK�g�
�"^���q���E+ 2w�<8WUqPf�XX�y'3��۠����[��ytf�������R����'Σ��&�����"���O���n��Z��������:�Ǎ�(D�P�ïD��>��1�f�E��+�P΀�KnVL��D���q��`�ㄭV�{����hQ�%��:�]�n�}b�Lr�O�ݘqۧ��Q<d:��u��o���'V�{rL��3_|#��WS����U~��U*��r��< �O6nj�+盠��E�'�,��=�$5<>��L��@3�'�r��lcl�^P�:I��� �n��y��� ��@�@����6D�U�o/�Ɏ�h��W�vg�+_��%�^6w�>�jX�^���LF�d)�8�~T���_��XG���o�F�R�7�$�Q��oHf�#�G\o	]Ɗ-Ռ��Cl���*MV�~ʪ���I.s�A�X��K��c�/��A�,(Yt�R컱�E�J'�7�HY3R�����)&�Jk&���-G	,�Q��Ys5W�'4hc�nf�K�T�v@���n�]��v�B����*�Z0�v���71����]F�#���#�۵Pǚ�'fR&c�@��5u>����r���x������sn4���c�PU5�l�����R"f�\��_��7mQ[W3"i�P�9�fy[�"qA|�q��O�'�Y�~�
Wh�VM��~�ڜȳ�~�: F+Fn�g��	n����e�q��(�G7H��
8'p��[����_SVAgǠ;?��WP]�*��D&��(҈�d�):��1���S����j���8��}a`��hoK��iL��"�g�,	KFj��-'��a��U8P�-�&��u�9���"'�3��H��7�����@�O��@���c���������	���zʼ�e=ѥ�1i)H�>������\�^���=�`��X�x>-.����9�6���m���+=y��H�F��?���s�|-t&�$����Z{Vk�)F@>�47̀�hK�_"Lh��+o0��g����w	�l��Vx�=L���w��P�mߕ�0�H��ƌ�cZ�qs�	&�8��$-ٔ��i�b�w"�?��O2���W�U�Tآ���Yl+�*��bHP:S�}p�o���H������j���-R�����%�2�3~ �{N?0v�&Qŗ� ��8-.�o��<;��r��=��#n�.qs��*G�(�lMh��=�%'RfQcO��i�F/���Pxq0Ϣ��̀�{����-�,���1����f��Q�3��#�9b�v�2*�x{s�&��A�4�Ҕ�0[�$���%>�:b`,\�+)
�����n��B� �,����ί/�5?BG�	�FCJ�X%�m~5�	i?����;ֻMP>�nAS�"�̊fU�~<�;G"'���l�C`����#<B�2X*�F��U��!%zxL�1�r��AN��6#�W���",��U5S��sQ��
�3J��vY�V����:3�\�O ���m3��V3����D����^����״A�/X����;5��(�6��a��>�<C3�R��k��q4`��U0B�[Q#�P��*��.���c�g��m^ v��f���Y�cR�o.��#��W�{� ���MVj��GM�b����~�Ԯ��N����Nd��$���O�%���3œV����6V�"](����*�Y��X��.��e�4���̋Gq�z��Y �wT:���>�x�I5��,�D+�.CUݒ�{�t�e���in����$����,<�LJܶ��Ț
�d��.���j����0�	��<����g�M��g��嗃��Л��]���);)�Kpc-��əC��p���-�|ݍuܥM�J�U��?H<�{Q2 ymkn�{J�J���1_�"w�w[��8�5ess�:�N�q����_員���I�0@��1��f�Z��m4�
`a-�̤tL�iֹ��H9�TW����E�^B� �ʩ	�|D#&�����E�R�7��_�Jy黣8��r�{pO�<� DH;{�a���DT�s��@�8�WϯPLhD��I.HyF����Vr�vCc�Z4�f��ZS��j�#������y����U���<�M�uX�(�Bw'�ƺdW������:�"�b���/�ݨS���F�'{�N`�p7���O'>���8����՟co$P�k,�D(N��5�k�(z�T�P.?r5g���Ɇ6߰Q܋q9��Ѳ,�	wGX#�޴����O�'�	2��lkwԄ���:n���D\םO�jFJ3+�2�	*d����z�x�	K�y����2p��|�ǅbBV��9;[	�7-63-�u����{p�cٚ����O��J�Um�r�����Y�O���9dx�?m��/N�0Eջ�}W�sH�_��Y� ���ɯ�M�s�:
R��y�h)���+�N�%��V~2��?Es�yH1�
��t���Dg
p)V����zoڮ�F#�	}���ޝ�%����+W�n(�q���9���c믯J"���v�!!�n`G|���E��f�*��oX��J�}�A���ن����🟂a��>>�嘲c���d�8Y !h�IG꧅zA��`��3�D}�)I��Ԉ ���$Xg�
�kn6�n�9�hL����i�r#A�ϟ��C�ǽ!@�	�������FA�9<OSE������%�S(�t&�oMX�f������ѱ�An�%��ur.>���(�u}�(~N�v�eBC����X|�	z�8R=�~S���=!�dN��� ��T�JS�(����u���ϖ�ؓl�/��� �VU�r��)��>���w��M�9���� ���< � �Q+{q���°�_)(J�Q��EIc� c2�)�n��Ƅ�V4��%V�ѽ(`���E�NM� o%����g��̃�e0y�j��.z�0Tq�R69����:��ʋj��x��2��j��Cq�P�8Q6D�Ț<��g=	�{u�/P�A��暻�������1� �5�њ�r�.�*�w̖�)!|g��:@�H�n�U�h��!�y:	�D�3�뷉~�AR��L����͘u�tq��q]��CR��)x��3��|�*x���٦��"Y~
!Z+T�Z�\x�3!;q�����>�~���PmNv��ed�5����7�K���U�tx_U�ڮ^�3x�5w������ccL)K���2��)��n��zU��no�����9�%P��$�zc�D��v�ҳL5#s^�����e"I��G�o�� �E-v��E�%Vm�2[޻�������^`���_2��S9ȒkVP�E,��E��V
V�zqu
�H�:޷Օ(���#��K�	0��U=�U�e�����U=�(����,����s��w�O�;�蚒�`(������XI���FG����i!���ʲ�C��MToE�K�E�����<�/�(}���;�,�3(�u:�V���L ��v�	A��m��B��:iXlS*Giʞ1��l2u���ށ�B�xb�0����%�$0��h��Q�;S�i�� IJOh� ����LF4�ϻ���\D���{FcL�Qc�r��J0���<�i ����ƌ�^�%C9��`�_b�+��:1kݏ(�U��!׹$�n���c���8=�O�;�sǫ`Ś�;�)+��批�QH쁃��~ӷ����U�s�`aAzVZ�P�����pt�p��5�-0�|�ǡ�Vl^[�~Ш�ԯ)�S+�_�dwU1�e¶�|==�������
K�OF�����q�{�om��sln�Z�b��e�d)�OB	��c�{�}�W.��h5!y�-�r���	r���I����nr��u���Q�T��_�y.��wlx��g�(Y�+�/-'@�:��߼�h@kON#����u�Vj��g#f���bi@5,!a?�O���ʕ��{��O�����2���4�4�/�0ɮ_��[��7jxN�L�=�iԇ}o4��a]$�Rr���[#�Jɜ�D/-�S����U�P�Ȣ�悭��n��^�~�YY���6~���jqI�E�;Jx�z�̔�dX
�=���2��P\$�����&���a^W��rxQ�=��&e���#��.ǜ�bCz�i�:5�B��xo�
���G������~C�,�r�Sx�[�b�<���w(�w)fj��65�DHg4M�l����N�iaU�[G�>k��~�C��94�yU,���*���9&ﳔ&�mYꞢ'��@X�^��0䈂9ڦ����3^tL����P囁�T�A��?�f��<��kԪUc�H(�51�n�;�a�����}�v\j:e�������[��x�wUڴ�+�R�VE/ħd�i
�p� k/Ζ#-�- �I�C��#ָ��L���nq|��Os>�l���M����p{F7:��o�+^���|��[��7.�3�/�F��g��p�S_����B�\�ʎ	J�(A�G�ֺ�z���\�#IռG����1�a��]�����i��lwq�a_֪��h�T��d;~P�ݧ�e2�'�In=G�$'�q2oW'5O>�c�Cv���)�ё�&&����Uk���XL�C '����LիC �8�^Ma.��V�Q� j�\U���Lo[�q�������"`pW��8@�|�&�#$rq� �;{6����GrDѹJ�h�70)��G�2�|���Z�9�#���`˶�w�%|G�' B����֑z4:|k��,�<C��qs����6a\ɝ@^��>��ѻxj4 $�:�+N*�����B�~�v?~�҅����|L�>X�G�Bc�w�hB:�qV��7�I�Qq�`���& ���=��t��e)���
CJb�qL���(tB��+��a�F�>f ����w��&g�ֿy��i<?8���o�����<r򿡏��H�&�*J^ �0ullYe)��[dY�Ħ�4qs�eo�w|[�$M$S��U������%#c�	$�V�5J'