��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_���Ч�;.��9wd�,�Ha�:Xx�
T�:�{�Z����U�kE�˾+ZM��Z��M;۪�7��_��.�t�)�\i��,[[�J�FT<���뜀�4�KZ�o*�8'r���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P-T�SDP�|�t*}1Z�h��Y��U���`)u\�*��
�V��m�[���g[/�x^�(�c���(@�<Htq$�9�� ����cVw��}��yz���%�٤o�����f)f�$6`��@A����t�SnP�h�7���� �k�N*��c��::�=�8�R��V$�)�U`������t,M�	������#�_m(+Ы��PO�@�y�eN�b�&4�tc�$�&�1���ƍ��B���JB{X�Q���i��ߚ3�Y�@q�$��F��0�k��{�#���q-�	��u�G�s�9>[1�H{K����|Xޔ����ϭ��课���&�jSP��3E0g�a��T�^Im���L�uD�,��.dڅ5����!)�*z���[{f0�g�1+n����H���D�%��p����zD�o���$N�[{(�wi��:�ذ1���Y��i�ѐ^�+ґ���uwy`��]�,y2)tH9߀����V[�&�,�Յ��t効'��2�����+/C���:�?Xf0�C�I���MAĸ��F1GG�杼]VȽ9���u3ud����U2��׀N{�3�j�L�Β��-���i2΋�W��P�GI�H(�l��Bgj,��4;�t
K�aㆦ	e�]���M/���^:��&$��x脀�*���r��)bȋ��k��� �#��=L�-���I7o�#�i첷�{�"�Z�_����ta���J���@SL]�t��~�t����Kݑ5�J����}߂ٓ}r-�3̮�n�뭬V������d������]���������']�d��X:�\If�'���{s��xJ�~u�滽���k�{5,�49�M��Sm*eeD�3�S�Vb_�ł��Ytu��v��)c�i��o���wh���+d�����y�?T��2D@�^*Z��Z.���f�
l��P� ��͸4n�L�Q�:Ciצ�E�M��<7o(j��e�����)lc��{��7D"|��jT�o�j�����\a[N���f�5ۮt����E��|��~,��3W��:�����2�V��~�<yK��������L:D��;[vP s�@�"$���Z��<�v��l��&%��}�'�"�$O���_���z=5������?.��_Z�u-Mf"�*�=!��J�Co��k߱e�{�`�����]H����{
���L9�H�x�$v�!>��n�i�O8lI�X��p"Q�@$�p�A����|�gk�[#�0qz��F�*(�$Ft&���D J�����y��6�<d�tX�T,�^`�� �s��vCOTaRp��8q5����@&p"s��̦<�T`0�We�<֍�X�������6�?����!�����+Y{��dR���Hx|&��Cgڸؖd�m�n�к����ep�g�I���j8�[���j2�x_�$��f������O�������Z	� �7zR�hݠ���̓�h�jX���gu�s�7/e����~�h
�������D�|S]�J���Ñ�x�bW*�(ߏ������}��S,ݖ<��{G��y���~��7�NW1��5Q8���˘.���'f5��oOW�0	�M�*]�T T�ɦ�bMT�-��q�ne����PQ���j5�s��V�>���0��-�w7��3���
�l[U��Իz�V�n���#JXe���l��BRW�tH���đ�z������nq���?(T���o��p�0÷e�&=�&����\P��Q���l�daM�:8��^?��1;�qc��9��0�W���hrzQ=��v�����"�{(�����4O����ּ
��b?�+]*���F�Q؛�gQ��[�e�;H~�kOb� ��Ix�/��k��񦩅,�=o��@��7�*���QET���<V�P|�@�T4s�-�C�?���A\�Ѿ�`�]���\[�^s���:�V;y��q�M왚es��t�Z��̯��ؒ)�}I?ٿ7�@R,r�+?��9�� qEhEWqm�����r!v��-�#�Y�������<�~5#Zn��A�"�Y�e����֘RLTс��y�|�S�'�a�I�px��)����e˓��H{y�Ŷ�
9�8�YVz5��6F���z�f���A��D%<3��z�.�(�0LO}3[�k������P&Xs�_�k�b��$!���7�ƫ�]�nG7>��j1٦wπj���q�"�A�ʬ�_��c���PjK4ݛ�����H(������OS��T�Dohc���oR8���ÿ�X�ՖH�6�#��R!�[����7	���-�5�Z#�՛K�i��#&R��y�L�d��|a�1���|�V.�w�-��x��F
�]�9�ȤW�uG5��Mf����$m��T�jy�g��BzY9-����g~��!������7�w��"�mIX���m��halI��>瘔�>�h�X�kƷ�xT����o<@�`3K����jE/������et,��`�����q��v�D�Ⱦ�@�8;dc���K���N�#�U��[.y��<hv��h8D<����r�,u��A������fNN��wW��!��ۉA� �K��	ZB;H)���ց������}�����̼��C�� �ƻ�K�	�*�0��)q�N�n@��V�]��B��SKJ2 Z~�͘�/9���)�6JX�y�����"M���$��sD��it�ВM�� h������`��ms�]oT��n;�BL�%5�N�7��Ew����4��$C��;գ �`3[��Z �-�d��d#��H�m���ZDbT�[IoPs���]��K|�HA�j
~< ��Y{Z���d��%�{�Y�x�9$�)�Ǣ���NٯS�+�4��=gp������Ȗ�W"�׽TD&=c��,`��f�Y��'S���6m���;�/�AX{-�i��t+��̙$�" ��ʬ�h�Q��aȠ��[g6�h��n�]U��fR�rK�п''���'�4��9��f q��t���5�\�&a#��&��cgm=&i���h�-�u��u�����p�P�b��/������v&\�g3�3~���WP����~������E���-��x=�D�O^��iel�4�]s��uz�Y�,�J�g�S��m#S�ޟ��΂�?E�D&{WAj\°�o�i�*���\Z��s�G�e���l�1ǃ}���Q`�ţ3a?��x�,�{-c��eO�~
�{��N�ĥ��\�I,yaQ�M'aE��d��ߗ���lytN��1�A���`2��Կ >���r1��z�p��'A3M��B
t^��A��~���#�*n3��.e=�:����tY�켹��iC70�?q;n;e�X�º(�����,�)r�Qs�XB��{�c��O�afpx�/-]A'�bX�|eKy�Ԇ����M�Sb�M��,��}]e��.�0���EP�x��oHFsd�z��+�b/�ҷڪ"�[r�:��f�Z�v&����%Τ[�m�����ӛ6`��.���w!6X�]T֟�y����Z�Y�ka�g!�s��$�h$�^���63���b@��	��jk����be����"7 M���¾s��g���i�}/����NO=������	��Ϙ���ۊ	���?@Q��#�t9W�-��h5���!v���n�0�̲y���O�e;l���i�_q &��c۞�x�U�*��S����T]�r�B
�-�?������J���N�|� 5��LK+�y��,?�w�7(ES,��J<�1�Cy�{��3ٳ�:*�N��ѵ�dJ#���##  آ��l)��[:Q�'�`�_�Xa��-R�1�LX����KGs���7Ѵ�$GU�u"7��u�v���:�s�K���SM^�Tm{;�[��E��g��f�6��}cud��ۡV#���<�ָi�M��Q	h%��t��<�:p��.����_oR���~���Ѱ�/�T���L�ER�/:�f�A,�8�F*٦�Uޖ��i7 0g���#
}p^A�σX�ԝ����\&�����4W�9�X�&�+A��WK ������?����}�����մ��  ����c����Ma��Ԕ�1V�r4g9nѯ�)�g%ߐ��u�ey�b�ñ�}���J�⠟���C�7N��la�\l	O״5"��EtE2Q�R���K� B���Jɛ�̱e �?�V(�%�'�
!8ب�$tB�oʊ�����}���ɢ6:�������}=�b�Z���j\D1p�9ߊ*���<��Ӟ�Uރ�1T}�`Z�T��.�:����u�o
_��l����)�JQs�{J`���Lu@HN�]�/����(e!xhj�M���dOG�=]x�K�ӧe��mv�L�=$�+b���r
2���������Sg�!�ut�V����<��=MNY]'�֭ C^��(�
 �,��&��B�ҏ^+�	J��P�qM[&��L\�%7�/"��I4�X��"�z�5DE�8[��xD���\|�l�v�Acĝ��נ�\v�1�v.8B]�rĂt�6H
��g�
v�g�l�!D����!2�᥁8�������\=�i0����鼂,���*��Z>;�G"�M���BQzMP���� �[j�Q�^9	�;��t������x�B�NqC�N�UiW����A�;f� �L���d�����K ����.�T�K���u�
\h��g(���X����w˕-�e�?Wq!eؙ8&��3��+��_�U-g��ļ���dˠ 0�\�'Q/EV�u	��	p�r��8��,>�S܉��:�`pv�0z���!l�6ŇL��kWbq�d�7�
�!��E'XEmS0��n� �^#�ؠ�ɂ�٣�KN��mc��sdI�A�������"һ7�
*�iĸN��̧�$�v{��� ���su�d1����A"�J����&�M��A|db�rh1�F��/+���Q�/Kt�#�l�PFͮ����}2K�'e�n���&�»w�JkѠk^��J���ҿ�6�H�g��#u���Ƿn���$(��e�}�`f�*R�ơM)f�hm�
2	�~^��t�:��u��*��r�"��:d�t���^7w��-����>=�Xqt1a¯�,�u����<� w� ���su�� ���($OM�V[�Z�ظ.A�e����Y�:�.�c%���P��wdx��#��!x�@U����˓�_�Gʚ9M�L��jj�.�� f��_R���Ź�]��8��t^� ���1�C&��4ɾaB�aY_�C�i-�Y����:FNS�Z�
���g��`�4��\,��Z89�ė��qK�?\�|������~QՋH	2����{v���_II`uQ#S&%���{�D�~�!�7�v��b��J_����ݩ������n�O�%�@�4b�6��k�j.j�͓�~�mb.4�jh&���B�nK����#�;@ke�0[���2��!4�;��
U20��R\-\�g;ˣ�O1r+�ً�?ۖ��ۮ{�p���L�1���"�8?�}'z?m:�CZ�wҪ�xG�؍Iy�<bz�A��=��Mjv߃:>]i�I\����v`��
�B�{MckzT>ا����|U�66d�AO}��� ջ�#>Hx�;�c��D�s�1Uo2��y҇L���&@W�X����l���i�@������<�%���ٵ]&��WY��S�I#��y,2��xNP���ҹ�3���t��`�-�/�N!�'V�Ә��һ�&�\jt�-�`���f�&���ΐ%���/���<8�g�#m���wF&���o�,���m@s*�#�Ӡ]��A1� �"͕Q�7K7��;9	j8I�6+����)�I�.�B����y�$4��z.|�>h��ƠW�]���\�y���yB�d5��q��e��$X��%�Ca��\�p_:�u	̢V�R'ݗ�Am``T=H�lt� 8�[�AtS��6��e�y�:��l$݆>�c�3��i8�K�mͻ��7N�2g�(�il_B�(��4pħ��s��P�hw�E[��8��/0'(^MS��By��l[f��i#����W��-$.�#2��u��F�O0<,�c��(�f|�+�ggߎ�o���;[rĶ�s"�j�DJwڶ$�ԑX���uD�g�F�)��/����,��׹�����5�0V�p*Qm��uSp�d�p��*���&mh��C��R�,>�N* 	i�� 1���r��s���/�3%B�b)�b1>ln9-�KM�S�2���z}�W��f$���f�Ma⟄mϓr���$��{>K�����e�q�|���B'�.gk.�W޽�W���J���'�V�ɗ�z��* �1�V�bqll��B���z3aB���Wl M.=a
���vs$�EA��Ť�h��k�#��S)�6���6���w��)�}X�;��ͪ�Ei��0�,�x���,eR����BhT����ӓ[�2n�=y/0�<��iYɦ��4��(��B��[q�>��4Ź��aT�����_\�Kx�*�>�K��)��Ӽ������:ee��Kz%����-�a�D�����NDf��v8U��AD1�6�8��49y�W�^�Èy_yW%����ﶎ������䩯���^�g��B�v3����~̜��C�$�㺒qO�QK����� HV(,�~�"�������`�@����F, &�I�1��0`?�Y�=�����b7~���6}�z�VZB�@�a�2��������2�����iɑ:�V�� �P[=.�N�@U�4+���).l��FD�k PF�'��c�'I��xD?"�:jL�tEUV���\��ieDټoF_�q���x��
R�i��[��#"��Fv��(�oc9��p�֘´0��'':��tצ�uw�J���㯈ډ�u�
^%��^m�T��:ǹ�O(�M��ʭ�m�~$.��;����]����Au�#��l����?p;���0�{�0�H�@mڷek��a`JH=bERƍ; ���ϵ��^��K�r=��6i��?��&�Wn�]$�Y�M~/���Z˓�ЊD�YN��xJ7�m4�oF�"M�Ș�F�E�
"�޽�w3ıʵ=1�g6��������(g��}F�&X6Z�,����?�%]�!d�|� ��R������2��r�%��p��
��ٳ���4�y��/�pi�Ty�j��$c�:�*�8��sO���^�M9�QM�Ϙ���b�����|a�-��
R���XFg���O���yfL��R�x:�qE��G@��rCX���r�eW�V�������%v���D��������Gpγ�~��N�ķ��ҡ�Oz�Ne���%�{�7�HO���إ�|�Y�rw�@荗%�����釕���eZ��0���ޥ����a�+�Z�OƠ2p�O��.�N�A�b��5*� a	V��4#Ghvg��?�j��
���.L
�9�!����"�L��	׻3R����uk]���oSLu�~��[��.��WD�ľ{|]\���>f������u�U�V� �w��S��QPM^V8z���I`�{��>�"��Ӏ�cg{էE6�P"<���Bd�{��hm�}�t�_ۋ������&vl�1+7�#_u�]���e��]&M��8���S9@���!�e�:�Cv>�]�X�g���E�'�~_y�U��E,�3���җ:C��[�������в/�KB �EH�SB�ј���&]��'���Ú��ڞ��`탯L�\2�Ͽ�,/Y�+�{�	���E�s�/����i��ҿ�Ԭ;G�����b'��499dZ�����
��{���s�p�l�$1��p�e�K��
'��.�ME*˓Mޕ|b���LT�s'���<���mu�D��������BW�p1��F��Ksx9�
v'�gF:�qv>��K��3	���$�W���/�����A�È�˘ƒ���.BҚ�<�� @�}�>v�t2�<#�_9�_c��V��Ņ�������d&�Q��r����d����f�N�j����A�T�h-}{Q{q�g���k��h$b�X���Z_��3��Àec�	>s�<~w�l���Y������T�k���I5?L$X��Um��گ7�(�M��vz�+��̧pH����.0���]][+׋�v��}H!��.��$�?;a_$WL������ɍ�^3�����@Z�e-�n�p���a�S���i�#?4Xv��rQ����L���k�;���y{��G�!|R�#p�dJ~��}'��m��WtE��%xYF,���.��d��^���⋆($�,Х�ş�Z�ףo����N���~|V�}cs/��E�tS�_�G㪎��ŵ�/�ak��GO�A�]��6��M��%����O�
�V�e�_�X=��S�,)���
��Ǫlx;�2��!�Z�K��Nވ��'��?�G�����B�	�,�N����i?5�.x�#�Ng�����Bh� �7���Ҍ��q�]�LT���yOKw�/.�㮈)�ᴅ�vV���8��6�4� ��{hU��h�c����-����y~�D73Fθ�AU �M*�Uootv.|Yn���b�Q�Q��<C؏�,>�^Ό��EBI��1�a���	WfW�(:<0غ������p���5�4k���G�~oS���zZ�	J�yRݭp��(M�E�������,Z��%��K�-��T��(��>{���'�_f-�a�2 #�>e�J���ܝ_���C���C�F�;6�vaܒ�Ȁ�c������e���τ�+��B�e�j�(�TI'���%1;�J�?��<�2��w����<�t]�杂<���e�>�k�f@������Yxqt��iI$��T���Lؾ�qv��N��U��l�軭i�>ϭt�G��n���J+6��|;�>�]�3ءZQ�IX/�K��^@��fGrt���3K	G)t��w:n]����?�ƒ��FS�1�e8<�5%T a�������ݣ2�sb��o�TT>�E;>6���E�,in�7Iq���{�<F�⌑�l��`z�Qº��h���K1y^r����ܯ@���8���I-|]Ս�5B/���ߧ��ˠ�q�dK���^�GwC Ҫ���	�Y�o7R�r��������PFy�+��g��i֍�3����"�-n+�F��@i��W�YWZm���;���%wL�V���"�ܼi�H��n�ц��גE���L���<1�Ц�l�ߘh"�G����$�(9bKzPˊ��9S�3��p�Nq��J �Uy���|�	���G�8�{=�Y�E�W�m��t#�U8��׵Di��Аյ�V�_�Fl�����pԫ�I���!����ǃ�2lTkS[&������E���sG.|M%�ۺ�".�+����;�ؼ���Ҵ�]��w�=
���	/� d�C��K�f���b8�{�R{�)Q^� �V�K�=lE���P U�l@}�kA��� F�ɏ���h�>�tumgw�ט�Be����dm�����ڛ��1H���,#	�?��%�� �c]��>���Ɂ��I��5�e�(�֟�����m�����l5���aj�i<�t5,'R�w��KŒ:x�-�P�_��+vܯT�U��Q�'i}�zl��	�B�N~	�MWSӻ�"�"�#΄��1U����+�Y+����0%�d���|"v�Ҧ��g��+�7T� ��Ñ[(e�i��NK�1���.�U�����ySz{Y�' T��I2.=�Y��N�y��5��|�{h�s�Ai�|/�r�B�妸��}К*��Z@i-}gD}�����g4��Չ�:��{�Ĵ��P���
���F�����'A�/>�%����K���|�W�/g���Ǐ�0��6������5����S�8��b(��'���aq�@K�a1�� �&v^�2�JrFіbǂ��=�K֞��N`����$��p�kr���}�M����a?�8�J]�v!Hp����
|�?��{0��eD�8�T�'�����.+ *&�Wd�d��eBFcs����w2�;����,a��G��80N�%��E`����e�;�#+�ݰsaj�x�<�!�zU�b߳� ɛEX��c�����=�\���YY|���w�E�:�p/3�ө�!�_t���y$�lF(ͬ!�'�j��)ܵ������1ܸ���2p�I�?A]�7v���ý�Ρ%[D�?��?'z�F�}�ʞ�ʳ��?�#B@�����!�4��7%�� ����P�_ֶ��+�(y-n�\o>�?@�����n"^�p����\�l��Π:��i��$(,�b*�,';[I��N�g.�YP�2��f� �u��4�X��,�{���?^�P�DS�^�p�B��+C[AT�+b���f�"��7����>����s����s���L&�Z�й���O�uk#��7�*�>S�qxhe1�Za^�����n�w����<�b69uVA�3c��^�wS�>�'e���\神��9T��V��]w�ނ�'��:gW�XXJ��������V����='7ʎݪ푅"e��]O0lTl�A���鴣�
(�l�;:�	+4q�e�����"���C�J~fz!d�6�h�L�ҋ��UG?��Ѓ ���r����Ztix���>E�yT>j
���O����MQh�Z�A�9��a�"./�����?&�
��7Y��H��������P������[����˷ZW����y�"�<��ZՀ�Ͼ՝>K�ם�҉9���8�s��@uW1�/,�t��8 @>�k�?����9&�r��x}�a��C7]z�7���DI-eo�Aҁ
�IZ�G��֎!z�x�'�SB�"����5�!�䤭p��&"�&��x܉��o�gQB��nѹ�^�c�Dd:#m�J{����Pm�#T4��Ŵ�y�}�'Ƅ��d�F�s�P�$մ��
�y����J��W�ꎅ�Y�8�Ƴ�=~y0il�d�`�mi|�Y`�� �����K�>�`�.��C��<��i�~�W��OG�HY͂B�_*&R;�`�cL��nU�}�2��ݼ�YX!z���B?�C��^4j�� �螠�/��vt;߿��/{�H�C������"�c�~��:����S�����M��e�aJ��:��s��>7�|7q­���W��GVC��g����;������O�AU��8�+��4������vE V��s�6d�O������<�K686WS����Pd#[���n�m�K@;KD<I�=����Ԍ%C3֓��J��T�ػʌy�msa+���O�!� Eo�B�;��tX�N�vK��jp7����fO�.���_���#$�p�&�kac�dG���g1\�&���Yp�JÌ&��tO���J�K�5�������~�1��9��]�����;�� '�U�{�KΣW�L�Q�WY�Kfw#�����)>�ɳ&N)��'O]����oaڮ�������=��B)�M�57ͼ���P��4r�6
.AV<{�C�����0��S;Ŝ]�@ċ��l;׳ܔ�Ǭ^��9%�g�����[ %8\�Aj�:>f�8�(�n�6 �� $��,�>��f��k+��1��Hx˛���Μ9}�߀�Cb��4��c�R��g��|U���=�Zu��d��R꫞���H.Ӎ��;��	�z�q�ۜmy��2^��XF�����C�%�SM�*�~�w��C��X|�3�M��3M�=G�R	��$~� <���7p�%�{0o��2guz���\���|�1O��@�^�W���0&������~;���.U��j����Kz���1���ib;��R��	��%��8K���]�X� �)�_��MQz#����ąDda���z|='D��v!H���dY�����%R���l��*1"�5�J	��#�"j�ק�-[b��GD}����9�*t�DW(�&~E�L�'�O��.����%�\�9�d�8�5��42�>
#q����
�h�[pg�v-ܝG���ܕg�Z�h/~%Ǣ,����Z`�Gt�mo���
KP�h6�<w���p�U��6�f�X��|eؔm�J͛_���m�{Z@V@TL�4��@v����n���2g�G�`�XZ�U�L�u*��k���|�����>q��e��r���>k�w�*���e|	�>�g�$�g�]H3�;B��fYԞ��/z��w�}���J�Q�q����юcW��"&ﵫ�ß�t,N�Յ�H��0�$����`����E��I}h�I:F�j��$ߎ�
�&�ț(R������<o�'_([d47��*Y����d@ng�(�3��
�b�����Ap�C������i��a���g������� �c32�^$2U��m& ��I�s�]��;��b)f���ȟQ��V�.��'�	�N�$&p>ɉؖ� hv�y-K"�ii�%��XJ �Kױ �k���B!�e ��.H=�ȁ�~&4J��>������`=0�뷈 o��W����?�T�Z��(�D�S���Ҳ�)�A�7��˒�������YܤimV\���"�q�J�'��}9RW�����q����@ �`��K9�3v}��i'W�ģţ���$�6�ݮ�aQ�Br[���A�����I��S��H���!!�!`��"gz/B��(��zUo�X��$�sLC}�N��z�z�U�GeK0�������r	W�x)L�c���A8�������k�El?F9{�.�c-�?Zg~$Ğ�8�g������7ג���׽Af�Im���:`����Jm��"`��*�~��|�G'/S�5�!�a%��6O���/]zT��裛ĸ�Gr�����"��X����k~D.J����UԬ�U@
̊t�pA�Ԣ;@��kFP���C<�{E�����j@�������`f_(�IP�j�]QHG�n�m3��P%)�I�1o�cQ�6�C��q���9�Q2�6��=�J����e2�T���9�Y�<���טة@@�FK�T�%��4�ZO4�?XT1�ce�CΖl���~�=����
7B��{u��5��鶘NSz�Y�����d�2�^S����t_����:Xu+�ev)%�_����7��h/����ٝ��\]H8�9SE�v�(=�/Vn������� ���l�T�����$��|��Q6�Ǻ_�$S�k�2UX{o�l���z%���Au� Ἶ��M��虼#���Ә6��d/��*X"�l�A�0��}�iYN��d�pޒ��e]+� TS#أ��Ӆ� ���BN� ����)~�[�I"��<#��]3Q�.s=q���@���*%So����9�����������-k��$��C�������A��s�zZ%| ͏�^�p��`���ƕ�o�� 	ɦ$cЬ��&����v�؎���g���Т�/�M���練��l$H��x�+�l�S�X�e��'Vig���=V|߷���}�������2q�{)����� c�e�m�`��E;y8�֥Ab����%��lh�oe����K����4��,��)@�o�;��e�iF��k�� ����<�6�n^b�pׅ�8:z{5l�Z��4J:7�=Sѵ4t
:�Ҝ�0��C���Idߚ��E��4�98��rs�������FL�k�yE��zL���t�D]�qE?4N��܃�Ʋ�j��3g�<�i�G�7 [��pj���³����(�����/�@:���yӠ�,�5�&G�¤K�A�#T����"��2.���U�UK���K�Ѻ_�������@`+�V���	��?�F�ߞ�g���B��5�	�K�;K?~L�*A¦ea�K��<l/x6�ɢi�.�.�f����݆�8@$S���?>���GE���j�����W�a	��jU��((�㿵��'i�܃V�S���P��L���M�\���xaJ��U�K���k�$�1�����)��G�:����Qv�t활�	Y~��1����^���|�B!���"�;�������	?��Ƿ�΀W�����fJ�Tm͌�3Pށ�7I�P����K��6u�x���t�f%&�R�K�q����Ъ��X��!X����Rdu�^�[^��q,�@v=�V������Ɣ�!�|�Ar��{���{��[̎����Og�7��5��<�xԱ�]�-6���>A��U5��^�RG!��$�u6����r>6k�����;�k�F�Yj���yW�/��ڧw��
p����h�=�4�1��d�lXF>��nԬ����;k�j�5���m�%�z� ���Jq^�d�u�u���)E�bJ�o_{�j8� th7J�e�I+��i`�.K�Њ� ��|��FD���(5�m�Y۱Q��S`�5�F�4�� ����%�ɡ2$ѓ'�gp��~,#KH.r��=h�L��$�V6���B&�sߧ���K�<a�[I�6�Ҡo����h^,�b&0>�ӏr�D�vc7D������y.��p��]7���]v^RM��?�I���Q&N%F���c�Vu�`f*���	�n�Ѣn���u��n�!�5~����{O�27r��Ug�C�gM8Q=?��t�B�up�|������Ѭ4�}�T�腖V��pV7���~���[Ň�WI*�7Y`��#M�'�B����'ͣm��r��k$�M�W��b��'ʢŞ�	�A	�R�]��۔~yP�b|�!u�m�� G��3��Dګo��-4��YuӢ��2/�� ��2�����M�W"�8
�^r�}B����l#a�\;_`����3U���1s�{C�M�D��xތ10������P9��#���pb&�� ����pf�K������AF��o`Ȼ@a K.T=�7�C�/���o��
ʮ��7�7D̨�_^E$�U;�Zs=�}�Co�Ҝ���z�o:�R������q�	��Z��Y�D
�WbM���f���q_a��q��H��K�eP��N�A3|L�����d�4.8��:�ߵ�FIy^�������b�KL��;?-DrD�,ӓ�I&щ���^�֪LE����8'�z�����hg�ؖ��]�R�f�}W�<��yU���}�B���Eb�w�B����{T16v�Y%�8K#�k�r�A I\���0ｵ����EX�OJ]Cuw=��Yx�ӂ`zDH��R��Km�����?���^�����4�����e����v;������/���5ث�^ t�h����ț��b ��P�I����3�l��̛B4$����a�ʕP�Ӛ�k��:��8��0���h�����b���׍�b��Y"ZE
/�_M6VK -�I�3DO;�c���Q�|��#̬V��n�QF��S��|��7�0��,T8N��O;�C���a2�d��+f7�o��"�}*/��Br	��ay:Q�~ƌ��k��d��A-�P�׎|�pTb�=�X���i�lQ}ޥ/���nDɂx�'�s�&F.�����B�9�%\��{��3E�6���3�,�hQXƴ�94���NgV��/�n��ϯ�n��~A;CtW~6U5x�	e���� U�e��4��H��#|���E�����f��@hi3gD�Y�GYmT��H�.����2*7�L7wY��Y�U�g�5���E"��`.����8)�7�Q�Gf 3oYUޙ�� 9��׃¼Ą���u9�c�h�r_���vԤ�i��z�'�Y����菕��Z/��G^r���&��ڑ�<}mQeM���~��|�m�̣��O��w�ǊM5�N��1�3�(r����qH����q[&�ݘ��>p�Gv|m�̘�~�'ޠD���H��SWoE7(���,���bb��I�:n!+��$�fs���rY�R��R�ђ)U��6\�Ay,ote��lX�,�.��
h��@0x1���np��?6R%���e�.��U@r\�q�:�k�6߼���|]B��b�h�L4�6U%o�dl��fR�Y��OΑ��.h�ć� y��Ӻֆ���e��n�,[K�~�x�HE�l�(��]��"���|�~�fx�'@��{諵]kݻ1(��P�26�j��ڔy��
���ϸ
W���,��߰���w�aR���<�c��dqf)�oɈ�{����9��T��Wu�J3�:]Y�S� ��"K���x�����i�.��UH;>��p���{�o�$_�p2�|Mť_�S�Lw��2gD�}�{8�@˷�fTE��[�B�2LM���Df��У�c�\}�9Z�]43���NI�q4�*^�%��h]��۲邮��\U��ZL��1/w�V�X*�5��rr�`����Yy8����\g!��/��v^�LB!�g��(Թ�9�+�W�Qg�6��~U�����'�ʥO�y'��ǋ�F���}	� @�M�R%��Gi��zH؆��L�3�n����󊏿�=�ɁK�m��������q]����aʦ���j���q5Z�f��J�f�� ե���Rk&]Y��i�fM1>�M�8���x|@������6QR�i�	�U�(c�<���"7�̬^�u`� ����'jWm��&hh��so���� �|�Ik�N֯i���V�y4|B�4G/�\��r|Q%-;�Hr餵�+��Yۡ�%U��YvN����i�e;�X�N��v�|���-�)�ioMĴF���o��W�l��P�^��<����x]�֐��	Qh/$I�@��#��
�I6����-�ۆ�1uZaա�������x�y�Cm���>�[�rH�3\Z�1�0	��#B`F��ѵ���b3�>㯐 ��0V����e�������a���(��(@kH�@�=�	�ba�gBr�z�6�q��H���vr�V��,��'Yу0�7��Eň��Y�tT~���J���J�+W��59�,RIU�!R��vQƦe �G��p�m�T�un��Z�"����o��vW�مAҋ��%���S|:�����O�Q3�W�
�'UU��aY};x�ώ�%%����^QTOQ������r,�҆8;<�R|y����kݎge�%ªz��4�.#���?-������!��N�y�R�đj	�����6��8�_^�kD����:�u��c?���4�HS�wdZ}����m8!�K�\����@�f��쎝��t�bE�������[m����I>�:�1�o��(L����uGw������6�"Tƀ�A�SM�?�c�{EG�z��{��ww�6lb��2�)#�"�}�#�w��dZ�<��6��
Ze���;���-���Q�z�v�>H�W�g�*6P<J1�V�:�ƹg7�h̄��S�OPB�S��x��+�ĉ3oTKJ�w���<;j��j��O9_���S���Zu�~����x[�YLiGz� � ^|�,gtC�rB/sP\�bqY�l���oj,);ު	iQ+v�S�]����я��_�Ӗ�1`ω� w_p��$Aj��!�F�]Y�~T�*8I$CۇR��6�.����Z��d�{L��(�O1���8׫�'S�ʨ���V��+W��Z�>)�����P�����m�*��90G؏��YcK����`��Q5�Jp�oI��Y�@� �Ʃz���ڋ�Ɂ�[�M�O�8}�V���<����e���c�Q9��0�7���e�	��x#�_��B!�S�v����$/'갖e��\f=P�K�����5��� ��;��\Q��� RZGm��+Sm�֑�
7��vh�tN5�8>���ꦎ�x5��BKb���9 �$��;���,V�ֈX{�d���U0d����m_���EȒ�,I�`OP�6'����;No�| �6@�0�l�3}������$�8k��4	a���/�h>��r��ťt��~/�I�x��/��I^qlp3���i#צ��C̼X|<X��Tэ} wN�Ǽ����ߤR���*���%J<��}u���i�0-7*��}o�(u�3[f7��]�5�Z/y�e=�)�$��*08WYP�䪷?�<�4�k�����x��ߊ�T�'�5�z��!lR�Z0_Wt�`&��P~�P�/��6���a��뛗v�/R���/�,g�������mU�������6|t7�5��/:wa^U.�q�zj��)�6��~�����V~�I��4s�g"XV�Tz�!iu��>�H�"'b��㾷o�]��zy�E5�K��|_��.�[Oc��l�\��5�]3�m��y��Zj��'�-�X9Z�/�}XJ� 1�J��(�={D�SY~�;ܡ�+ҬdB�[4Y�׽{^�g"�Ǔz�%7A����S�X'�`2<�)n�4�Ś�±�H<�c���}����ZO,�E��S~P�DO�a@1Դu��Q��9gJ�Y�k-
�t����(��p$r?�`�no`�IF� M	�����S��/�(�#�)�(H�1���v���'q�dЗH�5ث� S�ƙ�@�5Q�=�oS��c���p���a������9�𛝒I�`"�,H��簮c�RAs~/'͐y͗C+H��i��]����>��[�_��P��We��:xh9X;��M
<O�M:����b�M�� 0�y:_���$��3�U��&��4G^�N������k,&���C�r�,�{=�6I�G��ۂ ��|5»��Vͱ%�O��U��jZ�my��LI�P��q;7�k9���P�n��*ʏ����+I�CS�92cw��� �EY��l��4�|��g��5g��`b�w��e9��!�i,�����rl��혟/��mq���R��u+�'��~�����<9��kQ�jyΣd(,� .�^���O�}��8�^1r���6���7�X�i�w�W��ҕ��σGE �[�!GVc���6�С�� M��x�؏�Cl޴��=N7-��7)o�J����!�Q��<����50x��a��H#={���_�K�����{�_b����+y�'1y,H���H����俓�~�Kh�u��M�>��=�'F�$�(�}i��4]����i��䄢�j
��CC*\���xZ��:�z|T�X�! 6�o�3`�	xXD�6���r���/M�`Ɗ���|�׏�$v?pB�2_�B�Єm2�'���k��+�B[�Ѥ�/Р��K�Ad�;M�����3J�{���Cq�*�{�W�h�_j�R+��ܴ�:՚R	�v���ϷW
1~�����eϣ��sTv?Fϡ���ҙclE#,`��S��އ=�aN ]���������13���^S��q�����)���\�iU���f���B�@�������o�}}\�L�4W��P��5�R����!!|t���׳&H��0I)g�=/0:�'
w�������MC+L�̰چbl�Aw|lz�4;���C~��e3��wn����28
%G���@0̊��|���P:J�0�Ź�/&�� ϴ[}�J\��Ӷ��h�$}�e<y��v�,I���$�w�� �+��*3<YP�Hd�}�!˯ )�e������2��FW��~l�$������ć��5�|?����V��~�������jsL�����w~P	��Kd�K�!U�X��*���s������!�)`�e��	N��eF���l�`��pz�rS��Y�j��{�� ܻ�+x��ظ�w�����ML�³����}�W4] 9�r�2^�I�j4������Eޝ"��!��!;���B<a��w�$�t;�B�/�0zL�x���/%Paj�MN܊�?(���4V3�T���2����3��e��)��X�+��}���G'�Υ��<gA�Ϟ��l�x�ʮ�bt��7���U��P���"�=��/��?�8n�x�~*Q��ա]L���ɉ��ؘ��7Q��V�=�Q��]K����(�Y����(SY����j�!�S5x6���Fe�V��P,V��X�R)���؍�A���*���~���6�C����x-�6�f���P��?o(�b���W 	^j|ǆ�^%f��v��i��gV㷪HwK�X��	K���(T*Pq����H�6\�����N��6�LA�7q�v{g�@��
^���"D9�$��y��G=�C�ulB�h��M��cf���!g�ۦ��z_# *�(VG �Xu������r��ɒ�Q����[�����lZ�'�:�l�B�yW�:hb�A���9ݥHd��QO���V �6Ie#��i�.�Kl���e9LI;��c��ԫ�0܉���T��1ֻ����gQ�EN�oHQ������:|h�9op�P�F�� �Y�Ӥ�w��'N$�d�� ��
�o�䜖����&r���&9o}#�����7?�<aE&����e>�j���(�E���98��u��*��Xx�GC����� (��i�]E���C�*�}���{J	����d�(D��5B��)$�����Yy�UE$�v�R���l�B�~�LlZ�<馯h���G�,�x`� ����;�e�Am���|T��^gh&�Ǳd-:����[�L��보Ę���4���okpq��Ƭ������TS$@�-i^
L"��m(�I{&,�j����)�nW�3��Z�p���hZ�l ��R�0�ȨuaF:4�(��vk�mṣ[<yu&��ꈜU}�ᆓg����M;�]��bf䦤k�cxz|Iz��닶3����9�FǰB��]}��)ZVNR��t6��&I+D�o��g�y��=�v�>6�o���j����z.��=_/e{�إ��"ZA�ƿvsy�R�
�~W�5�A��q?���BO>eC����K��T��'�*�ۭiFz T�&��O�2v�N��ŽT�]�幻>���b��(QZ3�Y��4����wM���ݦ�L��H|Y*{����=?ģi}�Z�pI�s�hh�ݎ�;�=��U�M<�j�Y�9�iQ*����TSQ$ �Lq4ݻZ}�����Tֲo�ww��0s#G=�������;�O)/�k��Z��A`�c���F�4n�iN�ǰ+-�Y��&��j������P(�9�q�*G�K�'�-n�߾�7N�dFu�F��E>�x]����7&(Ī�?8���&8@P%�*��a!��{�M�6�l�8��Bl�0Mim.���g��Σ\!ݔ�Q�q/���4%���fO|V��d�ۗD��H/�C���Ӌ�vu����+ѐm{^H=���w��Z�Da{-�0N�tv7�F���O�zG�y�qo��¡9�ly
>�C�q���I%A_WA��3[	��kRFFg�J��?X��ٜ9n��!k���&��O��e�M��Pb▌4�"�hF\�s��h���>o�s�(���Gt*����	s����1�r�4��x�'XǨU���i }�1��l|X�5�-���T����IM�ʷGi�������ɁAA�{��wT5��Z�y�Dc���&SϥnX=�%������pAɫ�}�,��p��v�u�a��{�S�ۀ�R��y�C�_ww�'0i\�X�a��G?�y~�P��z��+�}�/���d�ƛt��LmP���Gm.C���@% ���\=�iX��
��Jޒ�@̂������;pm����E)2��9Nr3G�:��P<@|���+�Dx��u���:줬�ޙ*�W�t	�ԟ6��v&�������zv�3R�
�m����m�%��o�3�/�gl=��4���^Sq�u�x�ѶY��o�h%�J.��q4�����EL�����&����˚XH�E�������#lDbMq��l���=���t}\�k9���4��8͕�}Y��N)z7�+�x��}Xo3v )��a�:8�C��4�'Ǝė��b���5�_kWm����ܒ3�o���c
��I.���]:~��2D�q �I����C���ۧ�nc���}�D�T�[��H��WT#ѫ��/�2���� ��P?��#섍U�r����=X#��?Op�H�,lmF��֛%1h�)'M��W��ư�e劐&Is��d����.�R��>���6Hq��$��08hY�) ����W�7X|�$�1#ơ5m��Tj-�
��n�4�=d�h�D#QhZ��`�u�%B���%n��P������O�@6���3yo����.�t�m��^�>tm���m�ҝ��l�������H�$t�>�Gcq�����3�����wN��>�T����t?��].�ޛ/��P�����cP��xvA��l�T�#��Q4m�����~�kP�a�/������9K�퓺;�im�-�]�Z���29HX�
ak��V&F��"u+F��a����{��.�$	\Jn�[:�.�5p��g�Gˑ���t���XoQM�ͺi'�]�o�ΊtE2�o�;92A�i�?RFeo	Y ��V�����H0z�����=l� �n������E�Gd��$i�).�	�4�L�������o�=(��CW���рZO�-��RtT	��x�*���ts���@*i}k,��|$��;SD�l��Յ�Z&t3 �[#Ş�|^Jk�r7���bW������/A���O5M��9�,ޅP:5J<)�-D�`�~0v�_�az6O�
!�����y�?Z���o�U��ƫ�ũi܊eY�����͡��nT��+k�[T���jؗ���E����K��B��ib]p B7�R����F>Z���{s��8}��h�/���'�����6
�5��܆��w}w�9�qք1�%�bj���l}R�̪y���ո7w�1��[�-s��J�s���/Y^b����F�ޗ�]+Q��U��hvd�AIwM���pv��A�����*��|���2����K��T���������F&P]>w.kQ�@G�(j������A��D^��T\�6�rk2��1�m�~�`ȅ!��u<T�a�5�1uCd8�0HZ�G�=o� ��{���.��� <<��Y�����&�@;��q���:@�؅?�;��7�J8��BU�c3�z�"�Z�&ťd����=>�o�^Z�՗�e-|�Ҿ>��q5�(�Mm�H��^_�$^��m������2�͵ �ZU_�_\"�}v����Ŗ�3�݃�XR���ї�����WNԼ���Xa�8�B"����
�5E�
�^!v�Moܣ[?�WNE�+��TJd��Ҳ�
�ZB�)�o]9eB�����FZ�{0/|���t��ˊ�a0�W���XI���8]����Xa��n�<[�w^���f��d��gۣz��;ص�<E��l�2^�H2a��E<if��G(+�v�go��&c��<�j�  G�Q��Tf{�A]�"�f$�w�x�M�ET�c���	�rj��&��b9-B����G�����]���ZD(�>�X"F�F��Ǐ�[�F��ۘp=#�����k��.��,��H��AD�ں�/u�:�_�lĘ�>�3/Š�������+L
�Ri�8��Ս���e1�+5`m���������L(�KE���ƐUF��OQT�q�#<��,Mw���N(����Kp�� ҂��:��w	��
�N��Y�i��sWx��\�9K��/���+q�*�0�B�8�;xCD���e�͐�;j=>䫧]�'�]�_x�(�mvB��Q�N_�i���;�ThW����Dh�%㓒�\hl�-��L+ՠ;:\^9-�L�&/gd���{M�$�;�e��g!£)�s<Y�{�N˕bB	�����/d��Q����͹�� :�W�罩|D��)� g���dn6�|:���H/��8 ۘ���=(�-�g
��-��h���b��a�yWF\�>�����X/Y��/4�S!�a��O��5Z��#��(��M�_:�&D;�jf^[�Bt�y�
�'�BNو���ڭܳ��n/jl\���c��z�ۨ�?�i��D��ECh+����,%Ok.���y�U�$�,�������%�WB;�<��jј�&ƣ�I��@�n��%���F��^��҄?sq� ��zJ�{���P9�{k� T��L"��,�c/�s'�H�-{��������Թ�c�"�K'3�Z�!s��H�������S��ֈ�T͡۔���}����q�q�z�4K��-ɮ_�����FѰ��V����{
���n�r�-����Ց44���{�M�j)�
!��j���	(T�i�8Om�� C~�J��rԥ�q8�#��m@�ҖaF������ھ}l:K��1��)T��3A�h� �K�#;3/��J.E�W_�_s�����,F�_��}캺XkI� 	����U�O>8�GO�Ս#mDTz_7�Ew~`�b�Dϻ�uй�_�kQ���yO�Cfk*p��Ѥ���x�v�/*���:ɿ\��P0j���X�}w��/	)M�m�%L���v�=�i��|?��E�LF�߸g�ӵOdk}�. k}�"���M>���r�2�������-(B�״<����K���kܦ
�'���₊}kƙ�F�Ti�y >L3����-�8�xE�
�*}r�0�~��C~�����O��\7��8�/Eٟ|蘚�����:��½�Hq�*���&1�o�F���7nQ4$A4lt0���d�|>�>����G�WbV�{��WD��fJ�����8��hjP5HWȿ��A3v�] �#�݈,�-��tU)%�����>k��H��lٔ n�eϓFK�.���2<3�� 
ܼ�!�p�v��_����!���=ט���k�2���X{hcO�]��RU�����Q^yh�dyHP�bt<����'��o}=�F�s)Rͣ�I:$P5�1����D�n:l2��|>a��5R&��j�1/����;��u�rPu�߉�֛���:O�v����3���C�����R��~X�㸲h	���e�B�5F���~ـ�#�uKKY�f񹂸v�5�ǚ#��7P��=+�V��VF<Pk�l�y9�+cN�t���O-myg h�^Iw��Wj��ӼT��Vu��B� �X���L������@������BQu�V�`i�|m��X��S�������{9���/C��

F���,�V��̀>@���]O�򩦁%�W6W=X�>�_��C�����I��,�b���VS5NG����	�N�r�C�&���Tb�*��1��S���{�T����~=�A%��_1�͙_���~��i�ꀇZO{���NJ:�pY�d ��s�u����H�&�upfx�zM/�5�����ђ�@G���I���P��Q�ɫ+����>i"	�>q����w��_)�h�s�^���;p�	:�.�㳲�<�u?�b�$pɼ*;a<�MB񎤞��C����0V�o2��J�O�p�>�-�Ao�?m&�&�u�y�-t��M�%,
��?��Ƣ��-^1�ro��oIv���H�&,(���Л#�n��
�oQ��D��L�U�_-ſ�U`sFB~�[�f��ۿ���7�*NYTc�t�j��1�r�<pK��X)����PFt�T�/�������8 
��S_�Y}Ћfc	�7#=$��la�����-��F�mhf��Yg��8���H���5��8	��ԉlvS�\aq��9̏�>�a�cw��i�@%gL�C�Uc�f����
�`&�i�{S�$�Ӭj���\����ǁ�2��#jد���
�(���2,Yԡ���\>���2��M�EY_qTcs3��U%�,����Z��S����`���t!"u:�W�.�(���?|@e%o� |�U��ZK�o�rW�LX�ȑM�S��9�_����ef����#���U=������97n]��s��:�м�������(lb�ᔊO���Tې}���6�k�XHt���9-(��'���*�p�-�8	��_�[����xNH^\_�Q����!\9؊L���e�D	n8ʒM������~}!B�"����?�-H��(�����%���S0gT=�@�/�P+�J�oa�|W@�wh�v���mv,�*Ɍ���|kS{�)p0`3�� ~�3坉�}7��`�5[��J/P�k��� ����Z��,^i�[�Ȑ��#��|�����0��x@�j�ͼr���T����=��X��OfG{u�o?+��Q~�Y��,�b��E�	��	���uT|���;Q�o-����y��Y��6�%�5N� �N��t��)Y��{D2�tz+6�@��kkb�8q
e=����5�Z.)fg�$����a�CrV9e��/ǝG2�?Fb�q	�t�L��#	�0x����58����@	��4�֟}�|��8�ֈ�S��p���|e���~I�J�,>�̴uu�ϴ�v�;��NA�ׁ�S�Z��O����-���E!D�g�H�1ދz<#��8��E�0?)�HI���w�T���gp�e
	�*��7�р<��e��1_$僵(؈ԋ��F�����l�λ�MtX ��T�:Ze/k�W�]��2R��.3=���u$���kKNl��q�~�o��p��?���W4��>b�c#g��]qbL@�6ֽ�>��M���9���֕�I��D�������3��ä�ߤ�#���C[͎�݃�I�msnM����|�4~�����`~[�/��[Mhlk^,��b�y�f�J/3��5�(��e]L���`�N�fc1Tip}�pv)�v��������$�N�4��mg&��F���t�Q2?̨�4���Q�&��U�D�����u����aGsND�C�AF��Ň�'b�Z��#Ld���co�~��,z� ��^�:֯�����Ea|�SUE� X>g�a�>�����������$J�:{�TZ~�;��T��l���9��LY7ŧ�[�e;,����N2o���C�G�1�;zM�TI�G���h�]^S�xT˚�G./䈄�@��p��_"Ѳ�%f�*���lN�H�so�5��Xܻ�4������\�8}-X��L��~�t����t��
 �7� -i�#�^ ������	s�-Pb�����?�s�+'=��j� �aaL6T�����H(ޚ��Z�+%��S6}ϙ1~�&vB��~��Ev�i�?\�t�=S�/�[l��G[�m�������h������M�?��k�B8%�Oզ'�_�ـ'�8ןv�Db��Ex��n�}��bY��o�9 ��8q��P�?�r@��U�&���@5���f�sv蓍��D�m���vd��q�����$�C6U���*=Ȭ�s V���7�2�E?Ë�@�����0gj��w�\�U��Xö=�HJ�^��3��x�2�˨Mwŀd%�,�7�zι�!m�~p 
���K�g~m��IP�o����CG ~ڽ����pX�2rl�͞������m�8W�F2܀�A��w	cȸ��P���1
���۸�ˏ���^�)�_��Ǽ}[�2�����'�r����&i���i�WWm�3��?o"\a��t2r?�oL��bh��4�p����פֿ%8��<g�����S�v�<C���3|Z"����'ê&���%�4FI��\�?����7H�f��]�� �/{~C�o<V |�#����>Ōs|{'��^P#���,c�8j��_Q�K�{��}��������8�Ku5��R�.��5Mj���"���޾v�Cm;bG�6�I�Y���dd�{:y*{ǁ�� C�nN�L����ܜ��J-�Ե�3�Y2��T��͡R6��w٧/?��4}�<�]Ii��#n.Lr<X��=��Ut�!}ivc��7�G��}$ �2�M��:l*�1J��O���~����E럜�F��~��8Ȣ�:�-��/5�T�4��_�K�芟��bX�Ms`���������CiϪ�oK�.�HբP{hihX8i�>j����b�UԱ9��7�z���y���+g�p�gk>$e���Q4�� ����l�W12षҊ���	�Σ'��\�%)|5�Ra_�,���O+GU�{�*`�
�ن/R�u� �#	CL�8"�F@*&'S�#����i��ㅻELrX*�(�Qd�,��N��瞊;���߀�[.F��ϝe9l��iQ���� ��c�A�bGp�A�V��	Z&����R7~����&r�(�w@���N���rdg�$��X���p��i�^vg�y��T`N#
W�k�2+F���4]S��A���ԒY����P�Dv���˫yhWX�|!}R��Y=��6�+£�<,
������_�q�.�9���BSOy�S�d�
Q��;��[�#
�'���g:c����lkW����ћ�M�%��9ì j'�l����"=��3!��0q=o�H��x���5L�(�HcA��N�ˋJDeO�V���u�^��A���ϡ�<���w����|�w�����C	�����hp/�4�v�)s�s�~���B	nE�Hl�o=�FC� u!N�;��|'�S�G��3/A<��۳����G*�:����^����[_]������w*���aA� ���89�Rþ�a^���!�������O��v�����֩�������}_k�\V�����h+��-b�ߧC����/��~�5X�O����K
+/L:�ą�G"����m]���4��}�����!�MV�_����w�v��Rw�`Q�U��ml�3����)�*߳��q��.�ǻEo�ȋ�}�ED�9?�6�	Ⱄ,
��;��xu��q?�v���6ԭi7�P.�˜��ͼ��`(6D��%q��1�C�;�n�=`�-M������W���:��YM��s_�/�AC�_Qsw,�fx ��N���Z}^`� ��'`ϩ@��iQ����&���6�E���6�N&�8t��ߺb��R�'E�c��W�7���p lm�)V����b$�D�u����~@|ܨ�F���b�ľ�[2�ܯX_��d^�G�Ga�}ڐ�l��ߟV7�`�����˦f�(x����k��=���;�|S<bf)��c�E?��� ���Hfl6��M��>�]e�r�pҵ�Y=�YĆ$ۅ�����l�v���G�2Y,�� ,3��WX���{�X��O����2PJ[���A�h����>r���4_g��wl����!G��q���3/\*��q��z��n+o#@Q)lU�=E�w��d3�������banaE�x�}X��v����혴��9�
dB1,"R#�c7�gF�`pKDg�; V!�FK�_03v�����e������*-�/�s'6�i�L�s�@ve�h�S0��k܏��ٙ��X�E���K�o���Ssɛzu���>(����Jn��V�l��;~M�<i�4E��������Ls�0�]�� ��yB]�!�BB��q�z4F�v{/I��%WT�W������y�-���l�5�$S��YmnL�,�i�Dw�Z��۾؆�!��3.�@"YtaC�vLyi;��K�����g������_L*�}�����O&ގ��P؆�'�k��̂����KNw���(���Y���}'>��F�y�&�#�P��׶v���ڰXhB�Zo�j諊pg�� ��wxf=�߸�#U0�>�C�|� �A��|tv?���N��&�Xl{���H%˴[�Hǉk���1DO��]�.���^�
�䩷WW�=�77�}��7�&|��N�9
Q�-g��3�<�	�U��!��� ��`��Q~x�L>B��Z��TE�&�YK�;�B�Sa.G8-�v��ù��H�L�Y���"�" <���W|б��#��-��Xh�e�M�����T](�M�xr:�y��	�f~t�{z�,�8b`���c�:�ߛ���+��yRRN�w���f/��!�l���
l��������RY��C9$-�>�)�i6�ժ�mg�j쇭ؑ8V�]R,:�҃ps0^��Rܶ����)�J�_���-��p�A����yk�r�p����1���F�u*,>��
��c��Sp���J�8��]��%��9r��:s�ƛzO�+2T
C"�F�/��c[����Τ�l7�4�-D�6J)1Iʴ��*���0P����Rw�56���ܟ]�������h��u�s)Wy�-���}aݬ����YmyN�����D��y�
�{ ���p�O��^j�۠���K�tO��r�r�˒�Y�����R��������$X�.���$��Rt�������d8"�'/MbD�?���ú��[k���SE����1�>j�	��R�9}%�F
S!��+����ML<R��UQ�l974v-����~8�O�݂X"��\�Q����eG,?N��n�B��?1�Q��tm��{�1��eC�	�8>�+Y������<�D۾Ygl��6� p\�_͉ɲ����?�׵N��3L��B !e<�}�TD�ӽ/Q
i#{���ϙ�M/E�^���|$f�y��M#�<�����1�v2�«p����q�S2x<�(Q�mܚ7����&JI�S��Lj͞��u$�)X���:4RFl��n��ʄU�3�]>�1��LirS�o@w��c����柡��5�����������p�?��X�@�|���u��u!-�Wdd��|Axz��uUj�1�@;���E<��V*9��ؚ}Ϊ3҉
��xm&�a��@�S����?�?f����9|��D��0����. �lwT�[�+�D ������0K����~a砼AGq(�*8!&�g�������y���JV�jw8��U�$�<G��I�M������|��"��w��QE"������YPk#�=�����/�O��_��op���]�r���x=�C ��.j�V�#�4'#��&r��Ҩǵ�_}�-����|�P�s��B]J�n���������~K�Y�-�"5��Rm�Ϟ7�#� Td"?!�|�QW:w�r���	 }�+�����>�Ar�]������	dR�C��".��+2&��:�i���J��!*�n��`�*�:�#��$�M2�Sq�?^���q� ǿ���o���_�P}�~{��ѕ�qX)����Ї3�%�"�_�"}�7�V�n&��~B�A�~��1��r*7�/�P�ʸ�g#<l�}OպF#qF��v�H#P)��U!�k4J���
{-�=���v�R�˅L7�)I-El\�L�t�o���os�L�o��N�j	@��~�����sBn'~�ݬ��$ՃA��e�e�M�1�����m=�ÇZ�Qnj`���~��B�S�hϗ�a�A ����@�!��h�Q��� g�I��dl��~}��"�<���
��κ���j�uE�r��W�����T(�I�6DWQ���u�N����/H��=9�����|�������iF�P�U%�S[�d��5C��b1�f����M��U�]C�_2/����֪�c�A�T�q���ؓ}�U������V�>d}Ÿ�1�t�L�q��U9���JVK�`�5��a�<�ь��eȵ��[8\-����'c)�[V��u����`h+!(����|&���'/��1��V!sbs�lr�%&�p=#q�p�S)L/�_�li�#��u[�/w���/���@L0����M;��x��Q�'��C^���D�Ζ#wRI���}�`_� /Cy�D��0����i_�,T|�3+�1���I�&:q1�,�l�_h�t&_��0�{-��<OK\���Mnm�x���Knõ��:Q:<���EV�O��6�%��xn�ԀU��.�}Ap7,�A�E|���2.�Ï�Asoo0zؗ!AmbcP^�ӡ�$.J�2��%�wȻ]�[UgͮT��*c�RE���i��[�	����Cñr�|��>K�{�tQ R�g�q������^o�ڪ��e]ܡu�"d���4n�6���-@�E,Wͥ��:��)S�is}�Ap��+�=�ڗ| ХW�jp�ni��� +����#���u5Z�]߿�T>77��O������-pj�o4`� zgZ�{�d ōc��?�����(�2N�������h�o'��zL;�����(�[a����i�^Y/k����{�5���o�����C�����{C�l���Qq�-s-���:ݥ��\΋������1-iZ+_V�q�6Mv��Dن�Y�����Y��:�'`�e��a��sO\�%��h�s*V�g�N�Z��ek:dQ�!q=�rݥr���H�0�m���1�jۋ��ֲ�
�t��u)����|N�b*M-��e�I_io@|)�/7������ ýI�)�m�E[����&��1��Uz��Ͱ���ۼ5r�r��|#P��<���l��RPh�f�f"��;����y��sU�)��N܈��Ө}�Y�xX�W� ��B�f�Bٖ-�El��"K�/�N؝�K8�1��[@e�0)R0JtO"NXv���uh�zQ�@��yӞ]�#�:yQ��L>��� ��F
���S]U>�M �M���8����u�+��յSU�[��6�)��IW������ђd-WV��emT��!�d�i\�Px���M���w�N0�A�g@��/x��F��6���>��O�?���y]
+��}F>u-HՉq^P(�`:�Y��������\��e/��fy���}�	q���S]$��M�v砡u�����3i�Q�$�� �]�T�S��q�96z�X:���>n��f:��=Zİ��t��!�0�Ll��u�`���X��a�B�e�=�,���o������Qt_�B�� \˸�i�n��ǻ�T������%z|w�2�h�#���Ja{�niz�
дa��>����R/7(c�{�c�&�!��CI�am�Ğ���2B�n�>�?ܜ2qW�&�ERc-����ezBC	����$fӿ`�L\r�:��lڐ����4�C��R��́;,m�>�%�wH�x�S�H�]Ϳ]ـᏫ��*�h�L����D�b�S\y��+�^ŠoWY�2��n��V�g�>���hQ��җ�ޝa�)��ߏ��R�Z=x~����g�Lm����P�?�[(���~�Ƙ��n(��x��G�kW��&"��E�Ü�*i+�ԏ�c��)�c�1\�q`n�h�{I�4^Σ��i��h��*\T�n��z��oGotXs���m	�*���I��/����PT@[���ǆ����ob���#����7dA[WQ�Y5m�AEp�y%��V}+��Y���+BC!������ɶNn�U������qb�?�gQJ��L2uW�\�;%�����;4��w(�В" ����`�U�Ֆq�Ʋ��u�	x`˺@�Ǆ��`����\�-��?�)�n�R���i��Dt��5p�?8�0��?�V�R
xsui��q���Kb���
Џ�x�Wސ�܄�؆u�)<�ةZ[!�2�Z/] �A��\|hoD�]ߊ���R�)��`tY�#D�c_��G�!���;
�C��gjAS:�4��'"�����У��� �|,7r�ߺ��=*�-�p[83��)JTT\�pU4���m֬�+*T�F��-������4Y�TPRm���qz� $\�i�����U�l��@��f�󤹈��.z�Hw0x{맸�}\����JU�Π�O&���B8_8#��
CN;��<��3#j#��j|���+������b$E>�Ӄ;5\��w��`��w���x�� )�f���B'1�_v��s՚�0.w���}�E?e��,��yDq��ss�~_�$�N���҂�9��|:�M�z,P�t�D�O��V I�Ք�C�"wW{�DX�/K�T�2�hb	�G��m/A�}�9@4�{h�GdI9����gXh]7�x�u�	���)D�k�=�����ƣ@��W�q�o��`���*�pF=��,b���֥��f@��ʗ�(�׵n ��Z��~D�q����'�J�T��i:ɯ���:�+Dy�S����j��uUGj�Cfe`�F()(�6���<N=�o�=���Q��D��N��4����p�f�� ��\b��:U{��Y�t��5��.{��\��i�⛸5(j�s1��>VŢ������*�je���ҚQ����HA���nQ"���cq�C���GGN��v�����4Y�n*�qp���B^N�z����A5ò1իf��<�pW����N�x�|s�P�� ���a���)w	�y��˵���D��U"[!XjCA�>��K:���{�ˤn�@��&�Hc�����Ҵ5�i�vN��V�Ը>�6$�����t�{��[A�M��%T���_�D�/4	���:���2H�@@�.�&��JJ,&ǚz�����h�JL�b�C&��plF4�D<v�Б0����V��3�6sQ���'��vB�3�c��J�&:kvFsو۸juR�~-�}�!�T��Cm�a8���
:M��|7eKՍlU�g��z��_���+�t$	OEn����k��\R�4#{�A��1NK9a�dƻ�idV@G�@ET�yn��ϑ�ǲ��ه��w�:���+ny_�����H��G5x�N=��c`c��847����Ap�Qj`^Y��1�Z��޻���k�GϖQ-Eq\��d �I���Q]� �s;�ё�q��|���ţ/���?��Jr�ٽf��m�#��5��V��3�[�'�t�Z	0�8�;vHuy�5�����J@��l�m�_��q���Pς���G���篺Sr@��VD>?��5���|� ]�]ᙚzr��8�,n=Ze#�V��N+E�lƕ�yu�Ͼy�6��]c���"|V{�ьj�����1����2*�nb$C�^�G���2s�
@rVߟ���c�T�SL���[]԰��(ې�Tx4*�'��Tv��Df�9 1�35
2.���;v�����Y;D�	K�U����5�41�3�F�w{��()��e�yt���������gD��ϴ����&����&r`\�F�H"�;r+AJVR����L!�M�~f~En�]�"у���QC�>��+OL,�E��ͯWAXl��f7k��ŤO�-��������w���\yT�(0��H����/4�cZ�ɾ��Ǥa^���':����gA)ׯ���5�[�<1���oQRY��s���yW�n!ƒzZ�x�>�P��X�����Ѯ8��p�%d����D�S���0]��2��<�YM�����bNZL'Z4^LD=��!�%	�i���t5/?,F~�1G��(O�@z����`�p�p�m^g�%���1ޤ�:<&��I��l�'�1N>;�3VNv��P���cX`o��\��r�����n��p�4���Rr+��^ ���s�νZ�������c^�(u�Lg�h�ڵ�$��D�^��6;u���}��'�ni��k�S�]I.��7$H�oӂ1��J���)�V���e���ٱث�i��c���wj�&9QNB���U�S��)�Қ����� Gc3i6�~��s�!����!Rw�D��T)6�+_��S�<�[Y!�֦������"�uXуj�Fxh
qt��ߴm�v�>@�\����rk�T�]���p����j�i}�BY�@g�X��{�ƩԢr"�-����|�d
54oc�jtE��z�~�<ݐ�&i��zcϧ&�Ƚv��8@Nyɰ:x]R��״UY5[J���3��U�����Dk��2V?�� U2�t��a�D0�ߣŨ_?�lu�Q�Z~|p $�3�pq�/��gt.#��Ǿ�A���*Z�_�1��ߐ� ��N(S� �=�"du��'A<���A����A��r�Qq}%���6K�d��yx��2����	�d�8�c����l��ʵ�X���/�?$q�U�FV8Q�{��������Z�. ��D�iI�UCe�k��Fƃa�
';�U� '��)N�vU����[�,4�����i�YN8|�sa�s�P;%us��Y��� ,2��) G$�~�0uA��\J�y�h��V�X��Yߤ�~}뾇i9��:�������`�x��
��uN�O������C���d<��JAC^`lhS�\�ʑ���� ٧+���H3�r	~�o��P��mw�Fؒa�������ֿ.���5w��:�� ���od�m��,���k_��<CH��8� ��@���3�s�ýN�\"��7L-�Q�k��� �����U�[�X5��3�P}&��x[��<e��Z[h@���"9ƒB)�A'��6��ms=�$�Nc��xC���)D1|���j��'yy���~nŇ,9h��g�.���������$ n�>Wj�?����7q�d{Ɯ�P��lL�4G��녾�_ݡ���{dsw����ae�&h��ᴎ�dP����ND[�G��m�>���A�f�.�H{�o8�c�;	�P�cGxz�K?3���ĤeMf�#Jp��*�TN���:�!س[��x��.�����|*���n7�7(��`K�V�c��(�9� y��%��nA:p���gJ�!4^Z��*a������d��z*�<}~���
4Y����:��xV�p�����agւ������a�Xq��~<��z缚��%
U�)������<���#��ܚcV�\����;�n���$qC���_/?�Z�@�h:�#T��Ƅ�(#D��MB�:G[��9�B�}�
4��R�̈h�[�XAD�n�\�Ve6����5.TR��>1��bK~�q�*�3�������H���>���+{ǭ��a6�f
�#��;��,���ç�/�8��L���o�D��Y�G��ᰏ���9�;��B/P� ������W�ק�J�3������,��!P�*���e~��h��*��hy���kH
;����U���vsQ3a��B�W;��L��>>�V��H$���������dL
rG�����Z<�j;?S��$��d��\������&�y.��nV���ƨ[�N6�x�4T�G=u[	���~��\3��;8��HƇ ��EY�l�_>Oj�|�{����Z�t�Ym�5'��np^�<3�$����t���JE��c+)ߜ�^dr�n�J�Vg�I���m�a�_�k���M2�̟�I��Sw���mO�n/;4CT����|�e���V���c��SDq�|���la3�q�����r`3�d�G��C��^D�4��V����d�<�r��~pq<2�`�1�`��=���"I+��ں稣6�#=uzP⬩�QwR���yug V:U���,��3������VZ��g�R�
˖X,�\9m8�����b/���^�¢έ�_��Ӷ(@e�����Z�[� �X�XA`�Ȃ^����7�W(s3h*�����*VQh�#o͑�څ�O'!�ɪ?��+*���)���K�?�UO�'Ŀ_���p��{�<�"l�􌟡H �k0�����*pY&��mc�Χ�*�,�G��� �4�A��� �e��m�&�2��
�f*�ϥ01�Ѵ�L��YE�F�G�N����`{̬fl�@2�e����w̱^r�i����2(+r��P��eZ��+�Pau|�@Z�;T��0�;8;>64j�+fYζl
����:[ >)�LP��I��G��R~�5�iI��q=��-�KX�	�9E�v=H�����.��8ͻ&`�(oU\8��'��1(�/ݯ�9i�s���(
�2��v]z�-��+i\�C	��(���7Mu�XB�D�c�������@�9+�Ņ\:Q�HM�tPP��4Z�xF���Chհ������u�PO⩜��l��?��L����R�^U;��''����u_2v9�nOy]|j�&�|}1��xr!��zt�vb���O�zcK�s��/����1��VW;��=�4�FT���Z=�h���zM~n�;2c^�V��R��M��K���h
���9�Z��3Ҽb����.L�a�)H'��+rBk�̼��r�s_0�K��IY	��*�Vߊ�S��Em��9eS`e������\ғ�]�*���-�����1A���u��g��Hfp[)sj����Й��K������6&���{�D"Y(j��FV���&ld�pv6�����`|�O98�qL�
JA��s�Q���F�놨�P����϶��������p:If[^��1�+��<��Qg�6��QL^\�7�|��b��aI)����t*�gxAv�db�=(!:�RHrs�����7o�Ԇ�j_1t��l����n���P�T�ғ.U��_�����%���A�7�:�^>�;�mL�)�)N���,#G�W�l��� ��u`�a4N�z�kE=������>�	K� �q\����!�v�'�،�}���G?�KT��P��W�x[`�s))=
xO0�9�鷎�w{���>H�A�T;DE��	xN�gK)}h�ҧ����U�k:O]2N��H�a��W���y���g�{A����	
���!
������%�k�Ca& �D���4��b��-\�	\3pn����3C��jPO�$#������ ���H�iC��Ҷ�:T��Iӛe�2o�`������SJ�M��sS,ۊَUC�ߦX}L4pݳ%z~��'���F%٤����3�z���r����J�Љ�^5���Xdz`��2��i��f�:�T��(��D�d�el����	)�C <�؊9�&��"!�J!�:�'��q�Q���+��g�b7�9�@x�Al����'��H�#>WK�T�oIe�o�� �%�������n���|��N�W�I����B3S�����u9�4�e1���l^�V�IaK��֒͹�P�)� �EC��j
��{����,��ù(�^�!U�ل�[78�4�T;���r�9�@�;�����.�k�]0���d-�SW��z�Uf6�2��M�\Z�LU$�᙮3`U�O%AI���gN�^��B�d���p�ҧj���������]Y����sE�c
�<,g�n-&�d�D&BzF��(�7L�`!�p�F��^)��D�>Ǩ�6��]a�݀���
:�_]O����^o��Kٺ�v{���89�d!�h����x00��H���2�o����$��=����S)��ॉ!���E����3]���fx������|s@\�&�l����Q������lUPHD<�0::UiU���bGܘS'��;��Nja�N�	�rM�����}I,��ί�2�I��P��7��CW4dxlu�Oof�8��N�n�8���
�{&��4��|���!�Ƨ�aRC���9���ȚyH�Y5E
�6~{�2Sn3�Z�^-�+�#r�{<�&1������+�'����z���$�m�x	�F�VO����#�A�0kge�	q����p��9ø���"�9�d�~	p���ٔ���͗�Ѝ��m0u�!гiTIo|�06��
 ����^R6�m~�O��F�.��g��qo�����7�����M�w!E��骖�Y.� 2@���5���@�b�<�v W7y��EzJ�e^��:Z�4�M�P �lhP��E0��D@�"K���"��f"����8�W@3i�q�y���}6Ч�T�l�Q�3�c l��+lz��)�0���KH�F�qX��^ȋ�+��@����f	���ʫJ��׾F�����^
V���a]K���P���>D�RU��M�e[6Jрd�I������,�cp+��}����Ag��BW�(��w25��8m��FT<O��Bj��{.d���U_[�)���~A혰`d��mBN�%1{%d�7�'s2G��̆�1y�z��%3�wo��%�-U4���^*R�y�M�eu�1�����k͕��G��n�T����0�FS������!��fZ�8�$��+���.��{���r&�5Yci��P"�N_���0�8���_�� �Qmm1zOk��|&\�G���6\E����T� ���Y�UA�'$����;T�*U)u��?.G���l*}H==�쮎���Z�uݡ�ƿ+�r�ȝ�����u�.?!���c֪[�1�0��C7��H~O��K���0`�|F�\|A6�,eZ]Vq��l== �\k]�f�!�s_�[�s���FAvԄ��͛Eӣ�e{����z�e���cT�@Zam���M�V~��Un!4�)d��;���}I7H1�2τ`�T�w����o���d�+"��n��_	$�uu��>�47yFkD뎗.��ͬm�z�� Osx\�JN9��Y�Wdfg�\��O2����H���C.���󶖏YպZ�(DM����l�ژb���C��!��xC��R�C',M^�~A��B�\���1�m��9��X�Jˑ>f�o,9���Ի����U�^��K_�p�ʥTxK��ݍ��1_�����s��t�ǣ�0�⊹<�堝���>�8�����iC�Bۘa}E���Ŕ��&d�6�o��M�O�8��H]��Wv��[��������ޟ)U�_��Z܅�:��\B�c8.�^l3�(����p�H���,�` �H�e"̝o��}G�����G��L>��a*�~|�ǈW��V(v+k���غ�t�W�cI*}@�	j9��%\uNdk��<��ZO
i6�n0+�Zqd}N�+���p���|u�o2��yxV<^��ը���@N@�)�����bh�V �
�k����� �Q��p�JA<�����Aj6��΍sL9��9E��6 �iF�w��/io�ҿ��Q-Z����6~�3�4�����C"�,&�1�~��|�z��A`�{ ����`Vo���ub�r�CżU�����#���K��Ɣ��PRm	UVu���3n_]�8%����'"��
&̫|D���.?�Л�"a ez��R)��d![�zr+4��<�"��w���<3ˁ��WG+gVc���9w���G��_���/,YG/�f�/��l�EӃ��&��~FG��дF-��dUP�)�Rz?/k�gDs��QЧ��?{K��PM��`bz����4�C����4<]�m��ʌ���s���� I�!v5dBj���w�k���*p#k�?�<�+ە��p.߿q���T�֤f����2#����F�� �cuE"�e�	��△{�.-+���������'��'��Y�uI�%���)K�H=�z`���B�������Ua���*��y��	"$1�շ�~E%߻�ȸ�7#�nbsc�����������Z������<� ���1s��֭�8#1D�����gԯJ$hn�߈�����M��m+q4�8��Ζ/x7\�*���$k�����^06�MG��=G� ёր@,�u7����?	�t�>��ߋ���ǶhJ���
��,Ԡ�=��k�E4V�Ug#~�$9o���$��jz��nE��X�{��oFq;��L	���R�+����%�BC@N��^#�d_��q�K�9��`����U��G5�<�{ �c ���V|�T�2�����L[�EU�ɴ�aho��P~Hm��6�9C����ju������$�����A]eySkU"94G��H�)Z/÷�F�_����z{�F�x�¬s�3��%-��%O�=�7oj����N ���S����R5���ι��SDq��Tb7O�? 5�,���!Gc	C��	j��42�ҽN�������g}����$�c�c���zO��G�=��7�e�w^����	0�ø񂾉��q���1s�M�Z0AB=�5'c�lJ���d Ǡ_T��©�@mā��k��M�dw������$GG���⵸���!�D���p=y���=�z�ā�ndMʈ�]RM�#VN�r�Ғ3�*���>Nkp�O�`���< �ݚ��٫�/9��s�qfR��{Mo7�*IWXð�@����XZ�R���R~7�����^gy�U�H��T�F"�2�	�dXG��X�A�_;b�Kbk�l�(%8�#��Š�������4;U��G�O�0@;"C����	��5Dg�f�0t:�Ǖej66�������=k�!,u�KҢ&�����2%���#ar�͕#�Sn�0r߃��:���Lj���L��_�z3�O����J􅁱���U dę�,=]<���3�UJ�����? �v={4�`�e���8�#ᄱ�i2/{���*,��������by�s>�z�#�k��<���B�$]�WL���� ��Di��v`����r��k�l��#�.u���H�k={�b	J������������ǜP��g:���ꦒ�l,\��P���>���S��o�׿?�(�����ܡǲ�b(�C�i�$���x��b��l����E�Y�-E�p�"��ߥ�&��˷��qpΚ�9�6�\�Y|��|���	�k���Vv��7�Z})��da�b���WEN�j�Ʈ�$�s1�g���*{��4jMў�N������x�4qE���tFx�S����z����$�H�3��	�ڎ>�{U'��^h��M	i�%̚�u>Q��4$ �'�	 	p9�M׶�W�J3N�a�n���O(�m^_�"'�J}���󳗱��"����t%6H�0ݜ��ÌL&^N�Y����,a��km��`Ԟ�;�D�00d5��4�U�����p_ -�J�	�ς[�&�V}u�'O��fp�<�
�+u��1��E�q6�YZu��m��_��H�!���.<g�M�7V��aP��8���O���qQu��<(����O8^�H��>�A�{5�'m0�~Rr{��LX��R[l��#��eL�GZx*���o�+�ZW��S��eI��c�E��b�"�؝}����:�ܲ�M �l0J�~t�l���x��^Wy����sJ�X>Vo*As�N�T Y=5���i�*j���� �D+��U��9N��NI+a�ia�.<���K�x�ù��
���}6�ս)���i3�Q�Ũ�R�!m�IM��%��+��^��ބ����{|9��wa�%�d1�U����E7���a���a��q� �w�uW���hoי_Nխ��n�Fm����y]�x޺r���䜚�dF ?t��!{����/��9��V�Ӗ�̑-����p9��=᎞G�z����ϲ��VF	4I��V�P�����կ���Ľ_�eœ9n�`��	q����j-�: � M��HڥW�WFJ35a����8i�_m�=���?�F&�h�)��k��H�	����(B���N�g7#`��0b~$D�l�Y����zEX�:i�j�}>_�=���{H�P��+v��k(cχ��I��y��.
W�U>��TnSEw*�|V���|��N�,�~K4f�\�s.`1�J��+>]�f��RV�s0m�1ʘ*�'����?h\����F ���&.�U���s��6/UJ��i+�h{X�J��=����3A����7�x��K�#�h��54�c~ۗ8���������[�c��S�摜&���_%�g���7s���9����X}}K����Pf�� L"�RNw�tY�%���2�UWe�jT�۷B���b`F�q@�E�%8
~F�h����E��r��#�?�6��Z!��"O�H��)8�P�[TU7�"@	��w�8��;��t �֞w���B���N�U�B��R3�U�⛹U�=G� ��X�0H�9uq��m���:�0mh;fS�S�t�][]�{xx�rk����Z�݅�7]�m@.���忊�#�j�����Rw�ΞJS@8ƕ������Bx6)�'��dq����ɴaw/��,���E� ����!�ED��@��p�r�*�����!Eހ{=��hSZޜ��~�Є%��|�%����0��k�k��q*����f_\�%>M�-�<~߫��g9�u���~�齄�cB_cZ��OU�����N�A�"{�|��_O�W�¥&:���m����cg���MILc��E�
���#C_��˰�6�@��w��J�x�eA�%�� ~��2i�쭧�� :�b�o[�_���6 h8�=�ҭc��x����i��rC$��h ��.!��L��x*t�J�9��v>�R�yI�o�G��F�_@|*�9�7eS���H�F��3%${6�9^+S�	��V�uMw�RQ�[JY��ǦL:o�u�_���䡘O�#�j��&8謨��'��)8�\h����/@�R@���.dX��i��>"4���7ja������g�㤭pK��l��X�m���2@8B�t�F$7��1��Da�
Y��<%W����K�E��R�:�E֎�9�?�}�&ٮ�ˏBA��z�2�wwH�9�Nv�*5�%6=�t'2��폅���a���`���/�63�+Z^��5�'�Ɔ]��gFEW���> �%����<�ˑG2�2\i�و����^�0��U��!4���]0&�р���Μ��+�j��[�0w&��YE&�ln�)%�.v���uࠢ*b"�����cf�V�<�h|���uo'�R�^��6��z��Ӳ]�ފ.��Hi&�M��	���#U��R��!Vi%��U7�؛�G�!}|��U_����K��)�ˁ�v��L�rL~��\۴��_����fw5��֑C��*�5�Ü(���[3~��	�*��+�7 �p�,`�rW���4���'ta�8(�3��0��iG;�LSn�c.'����Pv��m��L.�	1��w��z�0���@��%N�t��>��?B�#�h�5bg5��Q(�N^̞���O�5|�l�?fh�Z�O�To|�M���~,�ʟ�4����KY嬣�ßh�/���i0�c-fa_yɉ�է�� �����"�uixM��Pv�5X���D��n�>����:��^��(�췓zK!���s�$��߫g��e���-H�D^Y�w��ĜF�K2�<�H��C͓����ܮ������b(�9���v�[jL�`�-]�K�M�=���
��a��e�I^��gj�μ�ǛjD�05p>�,'��?����\1������֦���dH���Z�U�ҍ+�*dp1#I��T^��q[3�=���S)i�]�6�T���}��OR&V��Z]����ha�ҡ�j]+t:A��oN#�z������JT$�(Fl��D�4��"�֧s�S��<�%�*yފә����$�rS��y٫-�qωS^y&U�Rn�� ��bA����p���+U|�ֆ%����)�cܘdn��
:��6�W�x�"�$T�t�z�F+�š��Ac">�����;��$���X[�C7��@�]Ի\q�!g�<�Mvr��O�y�#�����Z�n ���V7�	W\��Y��4��GN��~�t�P���P�v����Ȟ/�~ɠ�W)xNci��Yf�)Zϔg:Go)��	BC|�N'4z.���ޕwwfJ�\��#Df��,�����,d�x�N[}����{�P�I�$j�(&�g���u� 	��U&j�!�/��in�}�+�w_Se��w�Tk�j���jo���d�J����a���9^�YưC�fX�� ��	OCy-ͦ��ъ~7��+dl��Y:U��D@Ҭq�Y�v*L��Ռ�l?��Y5n�tqս�՘��sj<����i?�ln3lB��g!�0!e���%�f�˳؍ߕ�XS�i�P�:DP3�m��B r�JR�~�mMd���n�R��qU��.��� ��q�Sg����1ԣ�,�L�d�PuA <U5�_a������j���eV�Mjvtd�`�y3/ve���:� ���۫&�ŝ�ki�2�<JbmCs�$f���X{ēފ�9��Խ��Ŋ6�mm�2���BٝT��YE��3��
��|�q���nBN;�\h����,�ouh�g,�pY��F���"E�Jr�ү��ގ�H �7�J���*�L��s�t��<�&��kzGb?	�N�W��R(�6ˠ#�u�[�\�Z45�K7��<4�8?����9n�3
˿�	UK��h��~�+�:��it�Z6ƙ͋ɷ�zN�� �o?q;~�8{���H	,���=J��u��4Y?�*���3���M��9�+5��R<`��Jr�q4�N��x�CBv����y��i���������4����L����"AR����9�%h�t_v��rw�, �^�"��@�#���d?ᖑ�,�h��v��5D�d���� �+��b���9��B������Q8%�װ �z�.��4�t��(�ui��|^��p�{;9�S�+D��z�rI'CFN�f~�[��o�����C��*;���EC��XpW�����"�-47	r�<6����a��~����;�3��<�7�������0������Ө��	�@K_8c����M	J)
��-�c>�8&1"
1K�u!lX��~
��ơ~�CɎ�Yj^>W�P�K�=�j?�k$��ﭒ4q
.��]�g�}c��j%����>F��T1M�Q)�9��M2�����r�TI$ ��̒gn�u�/`�=[�l��x��N1�専{�{����g���E򅿣�91ߏ�H�h����W�`bP��'�����2��b;oߗ�����S��A\��b~n�����C�E��Tݣ�:���V�D|�nM9ǊbT��Sh422���2J�	�R����<�w<P�)l����v���u�p�H�]�2�@  �i��ǅ�V�fL#j^ދ�w oR��&��1N#u��t��W�xp�������ypWdf,�>�hf+`�d7-n�����(A�u`��[[)v�h�-�:�b�
-�������<�6@���A�i�h��t�%��ť�H��c!\2)�Ϲ�ߡ҄��}a��B��ﮣ�,�b]���zc�ޫj\F�G�N�3�eXO��<��f�-:�T[w	�����RsN��k� 4;����ځO�����m��+,~䠓FU�,2����-^�����8��^r	u�>�����d%�Z��h�w5�I�U��Hc|�?g����$N��!��Þ#�掸��.k��K�^�8�,����@u���;f���L��-��y�g>m����7��yX2-ӷz;Y�t��H�c)KnDF�~��}���y�}��>���ZYA����IR��8����Tg��j&JJQ4J2ȍ�$дKK	�n�:m2� /�.H�Y���9���������ω�J{8�2Iκm�81�sXU�R�}U���8�[/[	b��:�@�d��z�s�w�,⢳�U��r����ʅ��u�ْ�^� ��,����#�J4��PK�Vqq���	�*矬��ؾ�#�-�ؔe�
��C�hz�f �%Jr���fLY?�4}|b�T��.:!�7s��>��Y,��E��~ۊ�\y�jLP�z�c4k��?K��ϣ��C���A�Q��'+wMo͖�� ��I?b�D&P����\t������e�a�I��.$�>��Df@�^��� '౱Z#T�	�o�"'��n��4��%}�����Q��.�3|]���1������\�M/y7(@'A�rr1:�����G+��h����j1񣉁��ΧQ]�'R,�,Ģ��t�Z\��g�O��NP�؞�|[?}����}�>��i|N�m�%�>ηP��<�;��K]l�)�&q[�A�^O>��G�et�rb�>�&w�KYR5\XΦR=4)U��i�vRo 6�gi�9K��z�Qv.�Y�ޜ.����D��]��vQkѭ,~/u=�Z���ŝ��Q , �����Ҹǒ,:�*��V^uk<Wr-��F�Η�&�IUn���S.a�7�8j?�4h`+6�\&}��T(�0Q�i._W�p]�Rx	Hg1_c�_���m�~J���*�s$��MX"|�<��_��"iW�Ãq��t�쿙��=E�<�"d� ��Ge�*v|FY^6��܃�Q��gbg.9��4����J��_� j���>����k�f;�޹N��4�1ĺQ��x�d	>z���L�?ۂ����_�E�L]l��l�k;�0�<n8���Ag��Y��b�F�x/4�GSW�G��9pb:�ѳ6X�N�/&Z�U;�I���;�����~��q�$F_�靤p3[
LfĐ�J��_�vJr�Qʆ��oA?�༺q7�[mz���2O�^���E�g�uO�X�n� Ι��+�T�罄�*��Fd]����lW��j�/�I^9΍K~Ah�����-�|�}��16�,7|��mR��M�*����^�v3�f}2k�r{�:}�9�HQ�IM_���(���9E�e��SV!Crp��ұ�gv�8���y�����I�rr4ZP����vӦ�H��)Y�ͯwTcUT��)z�D��K�}TFU"��|#�B�y=(�x"�Zc�~)JA�6J��_3�f}��r_ޜмk�&R���.��]��1���#�|<+�O1����c]��D�0N��99T)�j��$�(YWұ(�Σ�Wz���.��%�pβ���Yn�iQn �/$xS��×�����^٠���+8�w���3��U�o�=R�����c�AL}&$%E��Q���PT���̒x��W��xc)��fOs�FI��;f�$O;�cB�����+��0��'����Tq�6���`�M���%f��ޓ��o��&J�)�.E%��^9:$2��٪B����E��1����"����O����M[H4_PZi+\��=].�bE���{8��+���+zP�+m,H�I4��dO x�����B�r.[���z�0V�?�2���Z���P`��1f!h6���P�O0�E�������LP�L(�d@s��$���'�Їu����,���
�MψBKZ�9.+XYp����Q�e0&������ߧ��������2�"���,���8,�čf%��J~}0�UQ�Zړ]��q�v#�FiBlKT�l
I����ԃE͚��J����m[na�X� c��X}v=���Ծ)�Q<^p�7����E�4
�����<��ӱ�L�Z�1��B$-GJ�'��LK�Ѝ�)��*�T��-��R$h��/�j}�:�
&�%n㦮X�R�K`='K����S�!C������Z�I��z�ْ�r��$�)�A��b��H���;{;���0�P���0�M�iw���s���Ɲ6� ���	m�f|\sVYr�]�5]WF�% 8�zu�|���#�%�Iw��kxHzv�iqj�ѐ�C�[��(cдe�AddU��'��^4��o�^��ڶ������qF>�v�H��K���ېp1}���:��F�y���J����V"2�mt��T���yum�\�A;uO�������'3^�a���:^w�g��
݈�����T��.�a��r��&�-��z\J��՞�I�dj-�����ч�=�h;����<��]M����26�ۘ�L�ٖ����@���@�l�7x���;H�ؒ�H=7ͅO����{��"���[-m,!�~�M!� {���Z9�����ek�7X���-ǫYU��V�l�=���,��]jM�G�z�[Y͊�j�}�.�ډ'j��y.;km�Q�,-��܌(3WnO%�q��(�#L�Q�K5Q*+���,���6��)��p��3[��h�B���[L�9'�lQ�F<!�e�K1�9u��o�
zM�r$�f�g+k&��_�� ���3�C���`�ݛ9�Q�瞸;/i�'��QKպ���&�Δt��)�~k,a��$2�6���p���d�ە�_ Sk�Yg���H���^���Lٱ8�4hI���iMg���,�m�\"���$"��\�A�ה��S�}��\ȳu���p���Ɇ`li�����- ��F|,�pqU�����񇶐^t�����(���r=�$���s�
�c�z��d��\%��:��m��(J)�כ�ܪ�U��2��_Nn�sBҗ?G,g,�U`9s̖����jˣ�it�˱q���;R/����N�3	w��X�̺{�1��7�^��;����� ���O����Eu$m�J�@Gp�W����{U"�`�e`Tx��ЧtwƩ�h���5{�����Ҩ�!�[x7?� q���,Z�:R���ڬ$w�W'[�:&3�[آ���j�) h~���}2Ajim4D>b��£X�09��1?y���^���S[���h��x(.���3c���3���]i��Ic��2ABj
�y�tkf���n S����C�us��RJ8��j�c���U�Yee�gXnci�Щ,��P��Ʊ=t:�P�Kƥu��:�d�/�Ӹ�BPN�;��Av�Ydx�	���0m�%�"�@��t�{4hȶ�о{t���W�$fX6��|�3�/�&�^	 i�Xtqh��]��t���Rnܝ�zAC	�<&|	�	�#���neVj�YŜ􈷊��ɣ0V��K��"����JU�����Z~�$:l�s���vP������;;�c8r�(��M��J+�u�c���%��$2QN��5�m9��s[P�:Y�Fj�	t�^W3+A'���U}�S�U�"���W_-Sa���*�zE8�d�v��f����P>~ԉp��:�Q��1?/�n���g��4�?:*m�i���K)*Z�87g ��"_ڗ:������8��A#l�c��L�5xx�"���ڔ/]�(L���]�jԭ��FSE]��h^�a}�ܛ������Ũ��L ����;j�PI,�B�3E�\0�Us7�ᄲ=�*�Y�T�`��c����#�]:�1eԦb)
��Vb��2�rA^$=b��eq�K�xIP����\+�((�u�Z�W���%E)��OgT{�t��I{c&Yz�≿D��QX��Ϩ^ݶ��ꟊ<Е_0
ÁD�3C~��q}�����v٨�!X`ȯ����謝]K�Re6�(a�]��pmYp<Pp��� ((u%VX@�rj���jiy��H�������-��[���ItH��>���n��N	����|9!��0cl�,1���Ї#^�<��r�5Ӹ��Z]�f|�:R�5c��xw8YJ�a�R"�j������@\3{����Cg
���n:m�'/l?�Wk�8�G7r�m�|
;�u�j�UY���V��؆����G���"�7n��ԓ^�O�m6�*�a���c�9���v2RF.�9��6AC�$�R��bFUv^+�q�1��0ar�@$ d�=kJG���:��;�.!Ѹ�az�z��cE�ף�kVd��V���խ?�,iY|>G����?��� >�ʒ)���X&�WYF�� 7�DV����C٠�|H�+F�����4��٬Yd��CHH��Pq;7�| �<���o[��Z�U�̗�.��?�r�x�9y��Ż4���Nwe2}��q�_�򃺢)"����!{"��A�0o��C#q|���DbF ���U�1㸶ܦx���I��z�󥎛9d"] �;e��_�v��K�^�8�?�����V�J��ɭ�9�2�Pٕ�
N�kU���zYM���צL��b�*�*���X2�_�=���ù@��:d��ǩ]]���bP3L�� o�vE�'�\&d+��@<r�hj���!z��S&݅C2�p�g�RN�{3�u�W�
�$?|r�{�L�rt�$�u�ы����ky؋\�*gU�n�W#/!�M;�!C�ȼ�B9a�<��n(H�`�9�bSK�`L���y��A�����u�%L�+�c�po8M@�D��9����fȨq%\)c�%�V"��6�L��)�W����(�X���F�>���,b%�
���x�g#�i1v�)7��ӊ���j>Ϫ�"r�V�4�0o�x(�~	�Ut9�:<զUxQNj��=��D�!Jә^�\m&l�*�%"���|jq�)�#ϯ��v\��\�"��4�>b�Y�4d���r36h/�3���ǰ�X]?��
S�Ir��{�q���ln�ȸ�^��"��J��Q�Q�v�6(�27|z�zNd<o�u�J:�e\If���'�E1�?�(C���F!N�R���7s���6�l�,���7'��P������L�*\cJꯒ/V�[Ǒ}5��D�ӵ��Y���Ƣ�_%�
�!�j��d�cY��A�Q��㕃_lڞq��5�n�7�\��Iǌ1�`�:z�-�9���,�Fo��������Ѩ�ot>����9R Wl� �d��{Ñ��|�����~��2�j�����Z*-	{����߇����q��mU�F�P}Ng��L�<&�4n�	�6��U�pY����EĲ�<Q�x��/;�Q�j �!��<:˚E5�,䷰����$-�K�̔��[���������;�@v�6�7��vB�y:gh�|\<h�����l�RZY(�+us���2�͖�N��yawQ,���ҟ0��~w{����1�J�ќO�C�.�����ۿC�'����o��Ƙ���Z^'My��K��׎ ���G8Lm#���ю�;�M
w�I�B����VJ1�p*�����[���M�J�:�����XdG@�3"W�</�$��tS�f�lx�E|u�}�{M���`i'ʢ��v+IFC�[?����	k�m L����\bB���٩��yD����B7�5_	�΂�6���Smt޾�LI�g�<$1/�c���`�ٚ�f��7N[�F����|D�����[�-��}!�f%���p��On/�����a[�B��m��?Ì�BqF19�S�����=��&W��I���m,x�Q�97�Lv0T�)�55Ʋ[+�1'��쑋#5�E��PW��$�׍矚�l��g�N�9�y𣙕��WW੏o0�
����ќ�"�����k�G�ަ��`;�^[�w�T0�ߎ����;/~�Bd<ŕ�>/&����{�|z�� w#�t2�<T�A�s����)<e;�%w����2K�0.�v߳Q�e�4��ːpo�He��1����!8v�HM*G֙��O!���$$@>�NM�������<�ؠ=R��7++�A�G!��t�a`d���BσNU琾�&H��X�s������:7ǳ�e�v�f�M���5��&��J�73k��R�	^F0�H9@Z�#Ҭ��%<2�T4�G3j��,TI� ��5�����
Pg�T��g��>9���u�]s�ax���G�#�:��"$W������q��!f��Vi޹Fk�W������~���&������"�$������1�<C�W�֜�N��:��%JԗO���z�U���NAT������:w�Y���ۙ
��FE�`~I޽n�Ԛ��d���x+`��<R�	)v�U�_j�)6B���ى�=p����QW�_��=�歫�߱��롲��NdZ Х,0f��2�	
+o� �� �GB8p3�;�2�8��s1�@���k6��%ދg��`cќI׽�ށ��S}-}��i����hU����ʆ�i&�ju7�d��Q��l�YE���8�	T�<��S�D6���#埙�r�t��U�V��ĩ'��F;z�s�(���{<j����ڏc4 �Pf�x3�J|�
Q��I*��2��9R�*(�n����Ͱ&�4k3Bz��`,i�(^Ej��Vpnj}L����f�����GQ�?_jR�?�;W��]�KU5'�/h(�|rWD^� Y�2��׆	W����9\�}�q���|O��l&2�����x�B�x�F�)^���I,���V��:�׶i�k*3�E@���)y����h$"Gx9��2�x$�I<�KQRF	�J��(�&����*��Z!�S��3&0�RC����I��$�����s�&p��K5�AN~�Ti��V��W�yV 6ze�݂Uı�&5�Cw1����1!0:�;�Բo�$��_rB�ȜR?f�H*�u�p�=憱;�,�!`��V�+t�[5s]jT�'	��J9s'��u\!�poJP��Q�,���g�9/����������. �߽��]���tC}lE`��!j��PR����V�qf��/ �6��a����s�p��~ח��;���h������+ ]4����>n����|�*6iZ�1_w��	�'�zu���ɀ��}�֮�&�ё9�_%|�C���u�*�5-ί? f(�l�d��Y�s���	�M �e>�\�}l ���,���p�p�>PCPN�	�1Z�7(�a��ĭv{���y
L�#H�ʪC�9W��Z�9�Q0b�q��T!%������2իߟ%�`�X-ᖭ�%݆� �HєV�P�cӃ�A3��67p�B�"�����>�^H%�_Dn.?.,�N����z���m���ً���/��?�q�\dl�#��b�U�y����[L�1��q�}RHPM̦}���ER� ���?]J/ėWX�@`ē͓�3S�fi�^�)Y$�y��S��t�x���]���z��:X*�DWƶ٣*��w�Һ��s7��a����'w-#�	�`ڛ��:��h�C���r*��ts{�R?74�o*��/=�\�\B�Ak��D���w����m��*QWf��4VH��4ƢPد)��P��`��2�?@5[�R��|���8+&�-MbI7CeY7���.�3zs��k+wx�TĬ�\�9H�'�ֆ����:'��T�擐z�����|g�~r_-��;թ�w�E9$]9�r3�8*�p�S�<�vl':������ z��2P��t/k�k�>��ڔ:Ki��P�!�×�%��{�p{�h��-*�:I�}��jC_���M�U��d��>?zF�;�R��y���(?�q�����lt��:ՐK_@�J��Iߟ����P��م��IC� ��<�L���F�U?�2i��#b���E����M�P'�j'v�*wM<}0#w�Ubr}�m�pe��c�uߧM9�vb�Y��gÿ��'�t��5Mo����P������jP��9�����$���� > ź���g�zhՄ�ࠬ�z2�*�þ+�Ƃ�9�uC
�?��Y���eug^W��M�{p��y Br�wO0�zX֓��Q؂R�V��q��W�B3�![�}�a�pi��K���I	��ٸ���{D`����$��OEX����Kh����р���#?�
�Z��ۭB���\������X�:��d�-�%n�8p�4aP�F�m�dPۗs;�qk4�����A��>���|�y�3e��E�~���s���I�U�1���f�c)����;H�.���1=�%��o�X���45`���	�� ��kݸ��7�_������ A���h=b��~T�r��t$F�����N��]��D;C���C���9���)�� ��pk����H�I+Ϗ?<O~�	��ʹ-s݅r5.��U��V��G�p�"wu�{?�O�l�Z���_������K�s�3��Ԃ��}���X���Y����<�8����P�b�WT뢇#�{$��U&|"���叹��S�{���z�����Ӹ������=[ygCa�!|%�_�}T	��'�����#��-x~�u�f��=�3�.���.L2o����NV��{��M/���P�A%�i,Wۮ�)`f��l� nw��Ma�����G�v��������Ш�J�aЪ� |e�<`�C��N1�_���a�e ZT�;֗_�|��ė9o�/� U�~�CW��E�虍��҄�P��� i_ �&6�D5���3\�+���[O[��?�Ѫ�:�
GGq��m��IU�*��Q�w+�nm��3}�XTj�1�OBa>UJW�ݴ}�5	������|'sQ�z;��lѲ�ژܧpeR����,d��_��@��|-b�T�)���)�Z����B/�<e��Lu4����	�[>�)��Mw��ٲ��7뢠��>��'�ȭ�7��<>h��ט������{�t�~*�O�;O����O���H�|V�I����$^ 0�{�s͹Ţ�V�:¡�cs��#BϾ�Mr��	�)���!|�����d.ӬL���s�R(cg�\�p'�Ũn�����K�p�w��#�lL/��@��*�ժ��1<�[�-#rmEڗ ���s�M0x��� �!�EW8O��ͬ"�����	W"�����H�Y��[$l�������.�k���L��� ʁ��ڔ�"��GS쵩�(�u��t�f�\.����@33&oi������{�U�lΐI��;��sˮi��Ȳ-D�W��e�U�}�^?������C_��-#3{��AK6a���̖���.��a[��'�`ٸ�0���vru>$��8EtXuo3R��~�P�)Of`�C���y�����J����=!��8{�^=�<TR`�x�뷁P�����Ih�0�#5�p��`%4[��Ƃ=̀���׹�=�����U<@���Fk�lW���aUD�6(�/�HWq�P�-��hm�e��J�T>IC^k��V�mt�2n��i[a��b��{�f�u��-ۃ�D#�������d�9J��κ<gjE+�u�"H���_%�c�~�7?C�N��*@�B���<�����^Ƽ��]��ܐa��i6�1/9�_�A�	�|��B��rȪb�&f?ԗ3�C�$�݂��'E�$,hX�0 ���r�3��B�	z�[sUi�_�ڶvK��8h2��%�V�V�)�L��R�l�r���Ҭ�0�H���TmZ�q1�݊k�~��od�@c�S�l�rX��E{(�2rG��oO�Aj2&,�WL	��@b\F�hN��dA�oNLe�i%Q�.��ﲊ��x�
.Ø���?�H�!���H�fE}��ju-�6b�[l�\�[{S��æ��\G:Ɯ�AV��"�R�l��X&�r����S?�Bz��P�w��ӽl
^^�9�9����J��9�6iz:��ua��d�t��9��5P�0r�л4V9@�� ����Lnd��sS��Ri9S��?rY1֊���]�������S춠A�����!�M�}ʪ��ј��$A�mT��f��?���m(:Dټ���j�������|7��L��Μӿ�R~q�����K�x�!�E�XL���u��5S�)����e�j,y�u�������䨄!N�b�EAiP��qfߨ�b�ܭ\�̖��S�Z�@	��1~�ŏ�+�Q�-��x�����9�+�g4<�!`�X����� h��L؛�m!�`B���
����(��s�������_��5|������l�[��N�;�W�c�`�C�Kٺ��mTP>oŔ�O* �����&�o��u}���#���ҍA_�.1���,�e�N��xW΄�^c���B>P>�e����_9R*�K���b:��]-.ef�|Nd^8���z4Z���nD�7���"��u��ု���k&a�F�_��ӷ�����:�z|i~6Re���Mu��_��������pJ�x�"Q��aޜ�c�b���M8	�.���(DC��_����Ϸ�Ԅ�����x̥Y�`Y����F��8���w1�Г�{�)�P>��H�؞��*�I���|�5�+P-�oT�<�ޓ����>��9����?�?�5v���z��#%�`#�ӑ��(L/��K�J�[	�6�g7!M�^���E�4�c��m�������w��]�I7�Œ=1!������V�cn����pޚo=�۔�Qd��}��4�(T迒+�(U)-��\&�e����[M)G�P��B@C���������
!�!G�L�3up,�p�$�i�5���2T����綻�:��(�ן��BQ��)!N�C���J���M��^��Kă�����n��7�B�+P��7+��P�W�m��^�V(4K�� �f���G�d~�Ar�{+v0?��Qϑ&� �4�m�H��8t�d�߉ms	�OdG��2��m���.t�E���Ο�*�)���t�{�&�6�T0�8�͕ީ�j���Q� jq�H))�d�߰��xR�, v���y)�@\'b&����s@��`ΙEl|l���T��2�T\�C��}���\Y�H/r��;��<���o�^�cd7n�#g�S)d�����s��	� 4�*��#I� ��ɼI�O� �%�&lr}O�%3X�!�a+	�$,�4KЋ���xOs�*��'T���fO����="پW�}�"�gщ c(���7�K���k�,���s�,�ԟ'�b>D��I����&�Z�٭������q,�N�Uj;Y��S�O��I�9�lNRf҅���׋I�'yB9 �2Ѥ�-3o��n5y.��|��I �8�'�GZjK��N�U��$7�؊� 9�}�j�Ͱ~�%�*7�tS;ޜx�(����!���Do����6�r)ؑ���:�0-��H�.Bk�@��lr�O�"g�rM�|�
�B1Xx���=���["�6�U	%8�����r�\��k�[V��꣥ p���ĵg��ډͬa�
*���K�b9I���E�{��*#���7�(�ᷯ�LP�~���k:ǚ&J=�:r�&�b���n&"4������0���>K7�/���j�?ֈD
^-J����;�.����L�D�П+o����g�ë�p�0)#ʜ����o��K.�K[_	A� ��%�U~n7X|�9�>4v���pE�tP������n��|�PГ=�d�|�>@�=t+qEw��d;��4�Se��`Y������O�vW���ߑL'�Ҏ��ZBp��b�fn!�s
3�aV8v��Y��Գ�3 t�
:˴%�������;Wu�Q^)n����~�{?�Ã�G�^�!���5���OD�����.9&&���<`Sʵ�h/�iP��Ǌ���k �Y���d���&ﰐu��B�$�*��fa���NŘ��n:A�?X5�G?I�^������	��չ�[�m�YX~�.�m�����������F�kڙqQ��V���o�f�R`u,S�\�$$�T���ʭl�C�k�`�趯�M�� Nɍ�S��
,[EY�gB:�2�`��a�l>���
���Dg�J�Y��������]�|4�'sԧ�,y<+?����M3� ��Kv��ZyC��^ҭ�;�T����~<^i�ӴX�ݮ�ء%�y/<;KQ�]<�1�6/�B�����n%����>��=	���yl����2��Y���gzK9�=/���9/����x�`�������/�eٰ�7�5ӟ�vMn���~�+!�o�=�GROt��C�s\�o�*�&�-�MX#<�����w�-��r%5,�R6H�"r���n"���X֪m����kVhu5ջ��	�㰝G8��>�@��u�l����w4?@������� }�g�!B��ķِ�=�ٗ�#�Q��"�J)w:b�`l=@�|9���� �>U�T*_�SEr�R�!c��R1dq�j��e�^T�`�9AG<���cK0�L^�����pie7�3S��9^�����u�m&#��[8��]MK�d5��G*���� �(u��sۺ,e-����3Ɍc	�ߜ���b-Fyw{]t��3�c��ђHs�T��XTZcvL�U���D�o����j,n�,,�t>�UG0Y��;m����њ
\^ڦ��?�뙹�Ƞ�b�H��|�:h�i%���tm�"���)�G1�h�t�,��۲��� �jM��%��<��W�1���]��F�W��Uv�E�ژR�Gb��]�Z�_U���/d߂#�LY[�U�i�ͩ\K@�U>�NK�6�̖G[)_q�sx�C�
��_%D�6?q����5�U˺.؝;O֘�=�b[ܜ�2s�j�6�g�9w�]�.���]Q�T�Ϻ��D1I�#�����g-����q���<&namLm��Z��ч��ۜ*�د��U���`^(�g�_cj����xD�t�c\�}�����I��湧E�Q��0�$��G�#��������56���9ΤbP�D�)%��=�H�������͊85��j�feV�:6�G+���{I"jol�{�Tw���˂�:y�>�T��L�,��	.�}H�q\�r_�O������Q� ���KX�d#�'�8��o�-����lY��H�qyn?-dwޖl�����<�_�Dp>�D���}$�?���B�Gh�E�ʯ�/e���@RۘxlR9��"�I2��*��[����Xkt�J�Y��V�T�#t(��G�i|Fl ��چ"�7���[�S2q��/1~q*��Vs���S���2!P0V��%=@9�5\R��6� <�'��  �$���k��r=�"`3�$+�^;ʼ��8XY%#��Յ�1�'�9CdK�W�ŧ�v�HF¸E�� ���A���`���hp�z�*P���c$yӧ�w���������Kd���K,������l��v�0loa�b�]ŉ��o掮D�@�-\13n\�w?sND���Iް�������t�1����1y��f��I�)�(]l��g�{94��2ܳ��v���F���4�oy�,�[�!�P���t4�[�0�Lmٹf|忲�T����l�Ǹc���B8��p�Ơ�^Ş4K��Z�ֲj
B ���<Jx;.���E��N}��S�"����_�{�W��7<J�$�o�LC�����{�a%q�Ʊ�3�%�-����d� �")^n�2O��\�Xa5t�SE�爾L��� q��f�C���,qNV���O{�v�$Z���l��w�m}�W�>m��y��b�OM��=� ,�E�&j�*�eB�Vx���:)�G�g�
/��s鋥�#^cںeL&�`8�چ�M��`W�p��Ӂ�N�*I��=rk�-T��ճ '��:� _6�n�pD(B)��Qs,�ca��
��3'�c�`mX��$�c̛/<iMO�������B5eX��u!��ѝ��y~��P�QEץh 14�b�C&0��n�ό��6X�2eK[.�Zu�o�Gʅ���I�1M�Bx{�<�/5�8u��z�VW����^�����w�x
X~a\Ғ�:*JW�RC��2/�YtC��4e�O���+��LrG�F��$�:�gKp�3;�I,u�'�ˤ��5��5��Tu��?9�O�!�`�|�=���j�ϯ��J��}��,)���Ԁ4H�=l�m�m�02d�]N+��A���[�K(��x�J3;�r����!�R]�:�[@�l�TveI� W<@i�}��l%��ܧр�,zDU:S]nS>��y-���6�l7t��]0�삚�)��w� ��KO�I0�Ie(T��hڻ؇�	�0kL���O��nS˲��#�5����ʒ�X0l�!5��^A5~Ǫ�=(�J�JnB�J1��E�����T�B�AI��F\��kid��4�a�>��P}��9��hC��h�j_ޤU���'*�n�F�T�_DA=�g�3��@��@羿��ײNEe?��X��%�}������G�M:��n�W��Z+�|{Wg�S����
J����X�!�p}��X��� �����	7���񨎹o����7e8��}0�YYo ��Hl4��	�Vr�e��/nU|��w׼�ėjE���h���)��N�L�%��>�ͪى%�����oT[�L9�&�U@(j*<��ȯ�Մ���}>��j������������Ĉk�x!��?�4�?%�������k6��v	۪B&�'�	7�4�w��s($�.`Q��v�����82g]-܆U��Rsgtx}i�1^�Mhx�;���U���qnO��$ӂ�{��g�܍܊x���9�β�_]�0�Z���0���¶���ǽ���J6�:v��A��ҝ̯I��X-x^'d\���+$|��J��lo]��z�f��
���@zZUS��T,�Ӂ�K��0w�_�z�ơ*�D@�n˷sb��L �
��d�A���uo����u�g��M����@�!k�^(���T�{�i@Q��.�D?�y��1�&���
��ҳ�d�Hʷ�ɖ�Lb�ɟv�m܃%���?1Y6x25m\05�����yV6�a��L�����[0�^~�g��Vm�#4��Y�3y�)a�I��YA�i#t�������A��_��+�TXo��?����;�6Hz4Ik�~!n��/�b�6�ƛrR�c�q��(�ܦ2���F��_��={M�����,9m7=�+��/w�.:N�l_ꁚ{5����V=�UË{Y���*��OH�A����]������6A����O�';��P�x�'�;bA�5�#aϘ�@�Ul}`�4� 9^v�l��9�͚��ao.�s��I�b����P�%�/x�w�G�`����(�t�j���HRS�}��ב�ʼ�ٕj��`�TdS5�&ς�;��j�O$��
Ǡ	Ȁ���A��c�D�H!�/+�Z�:pЩ�S1�	j#�4�`����编�(���͝4��8�_7��׈��V;R�3/�:I�~�dYTԋz�$����f�آEL�������c��
�ZE˪�? �v@PG��A:�M�e���.�1Mf���ՓkC�v�����V�:	�2��.��;�Z\����l�ʢ�َ\��,K������mA6�aw���0è~(�O�((��ꠖ����E��X��Һ��c�7sv�Xf���>��w�`������`&��hF7v���L;��Ѕ g�2�2�<���
a1��&�4n����8Xc(�v��坡	�� 4����=�C^��Q�n^�9i5)��c�^��UK�������#�Y�_<��X�ȳBR�,�aI�� jAO��j���UF�"t��M���[�*�x,Q%T��V��(k�~;bdU��*?nw���ՠ4)iMven8»��C�l$���,Ue�*�/�4���
FN�#H*̂}�h�U���{|�y�T`,r���������R�ru��[V�ݔ��海L�z�.����Ke������j}�L9镽��H�-�T��؈��䩛��W����[K�nPČT���Cq����b���Y;OmS���3ʞ����a\s�$.���7ʙ���S�>��#�����2c��ԉ?�~e���\l�A��a]ة�+���Y��T�n$��|8/\��er��&�b r�cS�^p�w$w�����)v{�5��_?�Q�C�#���Fw���F�唔���&�n��+�"�4s��J��h�ӆ�z`Y�Q��ۓ�Y���C���{���0x��]\�~!���
�?���I�Np��.a;��8hYc�b�.A^�Dy8bI����9��8t�]�D���x�#�4I����hK*�(+�F������U�½I��E�cW��E���!;�z��Śڻ��PmXO�%�N�Q7֑O|&}��z�3��j+I���$��,�p}����XS� ���(���nUNg��j��[�2�=�
~�C��4�yK����N�9-Z�+��1EN����ܯ��;��ً�y��4�y/�u�����R\���'5�vrrc��o՗&.�Y�y�y�~؂��3�!�}�ʺ���?J� ���3�J֊�^�54�ÄXƱ��pu���
nKz�'V�����9���\!���0+
[p<�D|S�~�	4m�_�T��*y��=�Y�TFAָ:~|h�������}�C)�a���� r܀�0�X)L-S�q�)�6�p�A�2�2�F=�ʘx��Ik�.G��(̺�x|:����L�����W'Nq
���zC)&�p�_�8����㴯N�E���!z8a��83�遇�O�:�O^5�H)�=����'0�'t@$B�Lp ��� ����lC_.wn�� X����[�ՂI�UU�
���}���Y���Nl5��[M�y�m�T\����������ߴ�&�;_�hW�k�3�_ħ�n\����qۇG7��|�Պ p3m�v�g�b����`<&:.�4x�������6�>N��s-}��J�D2;7s����������@9����hZ;��2��"�&�$sW��^�k�1�Y���\��`
��S`�"�MI�
T�<�`j4_�F���>lUGE=;���8��z<�%�h�7�=-
Dyj�u~{D�B>g®=^�vN�R.��ȃ�B�G�
$�jWձ�rŻ��F�`��*^�Gô��D����09	Pf<b�foI����9~E��؅v�	k����e;'��<��#���#{�p�7�#�]#/�F5dZV���XQώg+�q ^J�I틻�"LMvY>�7 ȸ�A�t�|�k� {�s��O.�{���ߑ枵��J�����E�>��*�����x͒�͡�l�	��K�"O� c��@u�u�˂:9s!�--�J.)IP� _@��#X��Ȉ�|��v^_b�e�t������?�29U����%D-R����+lU������uj�R���NHՑ,^�J d�;℺�����t���?�2⎗P��c(I�%��<��}�n���{gl�2ļ�2�m#���?|���_%�.���}��?�<҄��}�1S�w�m��j��W��؎W�N�\�NjH�﹭}G�`����^L���MF1��L�P���r![� q�����;VRg1�G�oo�[{�ח׽����C�4�"���5��n�J��j_��)����A���-�#&}�v/���+�Ǚ?���/lO�.�7;y��p  �0�ꘉҹ��M��}�ܑ�O��L�oLb�a���pE�;��a�f&�����7��g g�2{�y��.�3��F�l�v�&΀�ǃC� V�K����D�b��
է/ݞRf���[����wDt��l��K���k�x�%�7�؝߄��`�ݰ���eS/w@�}̗����-��8��BF�TV��'�L�Zx��8\>#�F�)����LTB������Q��tX�s�C1��C�U���EH�/��t1����+�;��ِJ�J�1��0�#�1�zg����Z�$8X�%Yb2���<�X=�V[hi �hb�b�LE����&�˥1��8|��ii��=�U�����;��E�����/�˜W|�A,�%���C-��IGh#黳�H�j*��"Ď���72ݺ���n�k���J�_6�������P�����bR/��_Fݱ|�s���������U�
ߨ<\�/���q1!�JLo���Q*7�1z���I�5,�7���_����&����
���-�	mlI���$�m�E4�vv�
�!���X��;��/�4�W����J���ȃ�"�G�Ԝ��7C����,
ј��p����-�toE��߼�I��|�G���-p�g�|ǘj�șk�s"d\`��V�m�S�XpL��	��W2�8�gk�>H�o`z�#��UU�N�Cy����#]���ª���*�{t��욢��^�i��B�n���;�j�(w���Ȱ���w�%��=^�'�LZq�����,�(O~��g�~W�C�c�8:m�g@$s�Ÿi�҅.f(��u�b?U�O�U ��J�'˦j�iI ̸H���i 8�%F�[L�'qr6[�J:k��-��*IQ*�/7�rg��� M�Å]�7�zKX�P+<���>���
bZ�W|���_r��M�ݢ���iǸ��;w(N�l���(x�B��ܣ��F�@yn�˖RSI���v5"�z�4&��W����Ҭ���Zs�uq�L������,/ܝ�َ˚�g���n�G��m�����<]�vI�~��j�9��A��2!f
��R6�W�&nF�T!��ғ�.��p�^��+��ڱ���_��6x���U�y{'�S�O���sK��u�{�eHQ��kX�ZLIWC[���x��(��� E���,,�lz§�6ywO1����[ăE9�Fll\&Hm�+{�6�Z�,c������DŽ�]�4
V1�چRS�<M�X��g��k�����gSҷt�tgqªm���߶�67��6�����tK?BXO��m+:���@�R�T���"�v6�����=|�;��R72�z;pi����!�t��C�Š�Q�'�����[�!K��S�S�����Mt� �d�Ys!��Vc_#���㪠�6��� �r�i�d�%*q�D������\��3^ub�#���`��tCNU&;�T��[�(r(?]�}�VWh���2V?�"ɒ$sU�ʿ:�wĘ��KS-)7�u���P
�g��;�%��nc�5��̿�����ῦ2����4�0b�T�,���������mj1�'�YF�n \8i�}�%\�K�_"��V�a��P�ޜ��f.���0�#$� ��7�jg�\sS_�-�6(E�aE���Df��
z՚H�a*a*�}
:± �/�Q6�Lz�9i"#�౔Vnn�rq��7�z�9y��T�K�h�۝��g2�3���/��S�!�y�Ko�j|��Ҁ��/#��p��N���C���B�2�/ni��c/��$.İA��*3i�5��}b�k�"qk�b��&F�k�~g�#���sW��fKV�%ߥ	���{׫LZ�PC����^:W�����;����ա-_lT{7N�N�65�Tb9�����w�9G,��e�r�� ,F1�#@@���"-�"�ek.R	Ϸ�8W�l�j�0��m�U�ߎ2���|7à��!���������f��G��u<�����?����j�143 $�QX�F��wV�d�1��g�׊l֜��Z_pջt�G�cQ\�^7��6����NG!o�e\��N_��pk�����}��ǐR�V-��t[_��vJ@lb����M#:.��eU{q���8ܝ�{�*�VBIC!�������=�XC:��T��q��XE�Z����2J\��\Wyĺ���2c����>��a�ws��P�� � �˨�';��*:\�������+턛����Q�r�t�s���R�?S��7��J�4Y��D_:C���'O͈���n���Rb��Jiz���)V\dǽFlSf]c�l�p|q�R"�3��"���tҒ@����&"����T��<�-D,'��Ql+`ƌ��K\��rʟ�_�2���� 
�>��^�������tHYzY�����"�`]Xf���W㡀C,J��&��E<x^��MQ9���@	-���u�ɽ#����*?G2�1���)��tc��+͌�S1!w����<)��)l�>ЊZj ������ >A��֦*�,	.��~����Q$���H���
9z�ʷ�5�Pg�n1u�"{��l��mޥِ%k=���ۂ��񌱈����q���F���EPKQ't5(T$"s�]�ۈ�V�8�f�٦�9��3}ӯ���k��������r�a�^�"�Z�j�b0 �Wd�EK'�9%r��s��*��\�#�v�1&���O64`ߨ�����3��r;\J�ķRM�:Q.�T��œ�O���-8[d�=��Qp�U)Ġ*"
��r�}zx�1F�a���<���[�KK�Zv�Q~p�&�sO$�д����'P=�Xi���7uM��%�o��~��G� �l���-&����k)�(R�I���MgSw1�@Ɖ�a��琏�M*����ɚ<����>g4n[|;Rr�IO���	ڸZ�V0.�tYj��d9��N_Q�U���e�ȩ61���gv��฻��/��?�{~f>��/2\�H�ً����o�����|�j��6H����s^�);�b��1���*�C���[�x�i��瑾=�[�h�舉��8�m]L�� u%y����-f����\M�' :/b�A�ݫg9�����OTڬ��5Q*�kU5�X�Hz��i���_�^�1��I?%�s�!a/�����{o�q�S��ǘo���4��b�C��m���mi,��E�Oϳ�Nr=�����,L � �]]�i3��b���ZW�T�J]%FEj�����
/�m�
�_��7F�� yV<X$�h�i���@�hܣ�5�͋���q3ǹ��DQ����MK������o5]DwVRP6+qN�	���������MU	Y#�T���6�Ȍ��?B�wuΠ|����Ǵ�����?�.W�2_����K�^��!j4t�i �'z�(@��q˓��y�fRC��CD�����SX����^�%�
t	n4��;�_�8�~�v����I�M��0�j����N�u�UU�ث2J���_���3��=�:VM��Vc:#�� i�jIm�rT+�	���Hϔf�z��:��'�
�T�z�����Eel�~�w7x����ДMo!9~r;2R��g�Uh��E\�!���ﳄ��!�3�p�U�}t�Nރ�؂<���7��vҊ���|��j�AT�E5�[�
B������p��I\�1�ׇ�]�OWs__��oZ&ްN�c��s�X����N���8���⮗�@:Al��5_�}d�����6ćN���p �r��Y�3��c�?g(��X�,x&d{��teb��k5;��e\$�Ԭ�_���4��L�E���E���S쩵��Z�I��*����K�4,5C��gi��1���Rd�;�DL!N�:�ܢ�:��>q�x�����!l6#c.�c��k�\4�B�E턼Spa�Ss�����_`m�-�ӟ��M�t��=�ʧ��7J/��@�a#P6��Mp�4�V@�'m���5�γ�\�Ӈ��aW��'_�u����ہo�	��'HAy��y�"�-���T�\��-�V�s咋a���
9!/-�^�7�>����r�l\�υq�π�/)��o�:6,R�#�p{�}��-���a������!���0����!'������v�a���M�6R9����q�V�u��sb�	��+ma�YY{�mw$���V������\&����J��hОg�{�J�oJ��Ǧ�6�ѭ~�?���X���1W��g�>
�<��d{�jI�Y�G4�A�}R�!{}MS�ᵗWn}#0ho��գX�i��&��A^s5*��?N��v�T5�����V�yՓ�6 ��{�B+��4yQܽ10�P��_���&� \�53��y�ߖ"dO,A�䭈�nc��=2���fL��S߸�5�Ǔ�;� %nfX)L��W����n��+t>A�Ɏ�y9徱wi��(�i	�b�E�9���EE\'ɥ�)N�厅B�`J�"��5�-�ýb�و�ƻ+�����z���0��J�A`�|)x��:��K��'z�&3EW��F�׍��j�@�0*ׇC���O�P���'%���zy��yT=��;`��g��a[MO�g:oή�ْ�uD�1��>]PgD�V^��_W2��ߐ` 4�ٳ�޲��^b�}+�ϧ���l�$�N>PZ �>$��B0JD���-Ek��iB��ǀs�rW�k��B��S�LhNs�I�`���nTt����g�v�D@�m?q���'��5��M��zf�pj��4��)=%��Lx�/�w"����xL�lB*�3مHđir�U�&<CS�-���DH��hqc�]����b��Z���������	S]��*�|��Y%ꚅ̝��)ٞ{��H�A�OJ[CӐfLHP`ٻ8��*6ҳJ�iA����G�G���L�Ar��ua��]����N^�(ߐm]���n;�?l��A8��K������U%jS��G��Dӡ��!E��[E�:f������)��a_3p�6����4<^,����U&�d8�`ݛ5:��N���s�2	���J���7�'-=�7��ͥ0\��6��p��TG��5Ŋ]����:����>2`s4-�1���8YϪD����z���������]L��#�к�_F�Dr�(tT�?$�i��-؃pMq$��"og�Dp��	�|�p���'��l�_�ы��r�nW��r���������m��n�w��Ӭj����d�<_b'KT���%��ͮt^����p-S�d���`\-Օ�Ab��?)��H�!X�߃�=������G������1��Q.�%����Sa��0gAqT儔ܴt�/�bJ�/f�F'fձ�գ�ʔ���_r5g��;�>i_o��d��H0*�m��Z!�Qm[={;�Y�����뛂�R-��5<�P���J�q�����3�VDmɔ��Ys�9�a�祿觟�l�������w�h�9�֒�C�:w!-�Xr�f���C�%���C�<P�8:��I����r�G<�]Jkt4�͕2B�Ŋ�ʳNX�O��D��RTD>[$��� 4F{��#O4��6�ȿ`�lu�bN�u)�pQ�}9!�p�]��f�.���("	����!�T�痈���.5�3����X�Q����XK�,,�QN��=!�	�T��h�0�����>9��KNU}Z�BH�Һ����eƅ�!��Ϯ��~�+m��JV!��K�Ѯ9���FWI.1֠�4�qsg�����(;mv=! �Ր$fM�=���0E���f��������m���'22S`��kmZ4�nA�ͭ��V�q�ܖ�Q�<`@l���S�[�3�����\�Q�\M4gЂA����"
�j���Ļw�c}s)i�9<G���n�nM=I��@W K?�M!��3C�cq�فQW��t=
�]�&��$\߯���[�F�Z�~�f���R/�ob���q��9!װu�	�(}��̰	�����܎��-��Y�����_�r_]��lB)	��0Z>)C���;�����5 Ƭy�>�G��23ذ8Q�G��w О�GR� �e�d:N3�s1Z��C!c��A��I���*�rp�*�џF>�
F���f���{$)v͏�H2����[d�|] $ߋ�?��X:YSC* ph�ò�P����|�> ����3k�3{4�SQ�T\��,Q��@[D`��+�df�;n5��a�ŕa ����������R��`�󿴿{����}�Ђ�;-���gl-��}���a�~�����BW��ِ�C$T����Y�����e$�A��[)����a����8S���.���	g�{)&��8bk�QA�p�0�p=��"'-���B�HE�H_���� 5;"�R��:X %�!Fi�̋��]ͽ���6�^����9�Wlg$kR��' ���i9x�(��_��x.��G��W����ӻ%�� ��i��m(P�������>r�
�/ S����d�j<�OV(�U����	(cר�+6T�0BKd�#��<�����}D����Xߺ��t�����	���:�i��ƦL5!Լ��Q!6��EE�7�)���(�T���z: v
TN~蝗D�����c�U�&�׎ ��� L'�sz��0��9n��R,�/bd?�2}6:!���Nw.�j��U�z�r��q(�
�HoF9��o��¥���H1UJ�p�C�gj������Z�W�f�B*x*��BΞo�`��Nu�B�sq���0���,�nvs	�:��c�!������ʕ�m1����ZKp3��HZ����w����9��Y[Nc��^uRz7 ��5sINp>|f�J�M�4��Y�h� ���R���j�I� ΂�AӘО�R~�c�0�o���;lc�-��GU��9�j������}5���O��F��`��כ�g���IYڒAĊ� eY�~��a����"����A�_�so�g����Ql�񿇿���(�#��;�nw�ё�=��F^=j���{/�F?�ov�b@��������Im��%DC��X�;�H���ut.�[m�{�=���U����8&x��yyF4��f�á��z��X�Fݖ,]g�=�G�H�����Df�F��,j�<	��j.��)��h�H��P�N�6���dz��v)�,���~:��pXۥ5_�)��E���%����	q"\�'���̥�}t��:B(�)�U��w<o3;�Şf����q�#˹/�U�+�v�Y��\4.9�5�����ua���K���L��/�{I�#b��+d���.kId�#/O�0�<p�'���`�(pA�t~�C%Tӏ����Y��m/��́�P?�ohd���TfL+oJJ�j%TR�Q�I�����~#q��O��s����5�Х��Y�f=�
�m���3ZxY��-\�%��*�����c���p�g���1�Ͳ�o ۓ���J���mZ(.�� �cP�d{P��\ڸ!���8��e֖����3₶��������FW�%��b�g�fK�|DFu�d��\;�-����&˴#.��p�2���O��m̘�O�7�!+_fs��x�B=��w����,��=>}�4�����VR6�f�0�R��,e��E�P�9��>&�x���:g�9��A�G`
��V\&��6�@@���k��.]�ET�.��p���e)f,�\oy�*:o��Vb0�U�mO�yI4ϔ�&�Q����L~��o�E��5Ό�Pӯ��'�UD�����#���Q~���x���S��ه�ǭ� �<����n�(;�]!�0���y;��Ok�C��-�v��-���9<MF�[l��*4�9�/�$���R�ꐬY��y�Fz��-�ns>L�fIp�y�"���iS'1����CBH
��A?�	y]�D�i�"�vF�x���������($�v>ʂv�<�Y��t[>��d�F��Y�9�A�%���=~	R�Lk�������Q�-_I���3���ب�ФJcكO��l�â�u�{�E���a����Ѓ��� ��1�Q<��$R 
� �8���7t����
�,R�/G�a"�n{2�-���Cy�����:�&��j�w�����G��2Dj�<Ƴ�ߣ��HP�]��g�':�`k����7��k�XA9�8�G��K%܅j����G�����y��]|�=��vdJ�}�87�R<�F�(�h�!��w�w][�㸸7+���t��\�L�U�f�1CՁ�n�W�?~�G�d�2b��������`d���]��q��R�KY����1*���2l�(�47���2g@ԇ�����EG�D����%��-߃�����p�(�����H��eFSZ�^���]�\@��. ���� ��GצS�u@�s�U>� ԇ�Q���"qo���&�ӧ�uK��{��5]����0+T��� e��-wO\�������MK�~��iq=��w�b�����h���<���O4�m�%e��Ϧ��2/5G?H��f8�ńè<�Yn�L>��"Y]q��}�M�.��}�pX�����.����qg%�������"�2t,�� �zd��`@<�ڱ~1�ѐ��n~8�U�q5q�ь�IYC�Yy�W������[�ȕ|a9:�mPb�t'�D/�M���vL���x���%��؉	ީ��Y��lk��&�~�aNG7����q�nB��ސ��u��eJ8��<bQ!��8��E{倡U��#+C���Q�Z�n>��}]W�R
$B�.�Ub�x��C�吢�zy{ˑ��
�Dʌ>wi&V�Z :o���Ǚ�ir���ņߖ�m��P�j����uvsY�Xd�d���$T�s�ȑ��C��`�ߤK9���K9"0�@J��k�e�nh��&�j�#A�J�Z�p	Μ!(I�u�΄:����pO�s��o�~�ڶ�Ij�N8�b�͡�r���HM9Y��Ƚl��W?��{�~�Ug餍���w���,��8��0�i/^��4�7+c��xĹ{NF0��;����,�R�q��Ʈ��
��t�b&�͞	vx��q�F�)]qP}/f�ua�t�;0����ix��f�h p#Kxg�	�oe\w��^<�a��D�)�p���8`�c'����^���B`����ڏ�ݧ�(C��)[��6U�t�=�Kw�0vqc���ݙ��4��7��LD�r\��U�M��$6�2�u<�'o8����v�C��$��z7W�����wy4;�ֳ҇�Ð�:�as��D���[�����}��Z?�A��M/
lσi�1)^�!��	�F���������c�'����f���h��x��՜�X0�7�$��ıw�J(�M�Ȥ3VY�Vx;��?�Ѫ�?�ֹgh�7M?�`'������Őf��� N~���3{;�Yx��j&�@h+K��a�{`]o���ø��ՠ��d@P]x9#��������ϵ��*ĥJ0�dY7�&�f�AЅ�Èq�;+,�t�K:ςp�#�������^04�C�(4���%Ǉ#a���ŗ]��>�I���]'�I���?�˽=�:PY����S2��n�����W3P�x�T?����q|���TԜ�
M"I����I(r1�p��?q��~�"Z���2]}��	mԶ�{5�5a�_g�@���kx�Qz�
��<9w�=-�����H�Kv,�O�k��p�PEв7C�o����������EL���=ׅ#h���&�G�h�˯3{����P[��p�l���5�L$��Ϟ�h|�5�#���S�*?���\�� r�O�"~��֝b�R�I�v ��"���(�PauR$ʹ�Fΐ���8(�����A��<^-_��-ı��?�� �!ꢁ�q!x��J���㾐R��z�/y����S����O9�1֯~g����F��:�H�����H� �8�W�i�R&�챚M��Ey"Q�	f�=OYh7�0�[FLS���q���lHx�TA�T�u>n��t	�a�~������/��(��YZ�E4-�b�x�"���W��d�Z��i��ZQe�y!k��ȓ]x��s�Z`��	����e��4�&���
���C�ۢ����~�yU^-��6gn�ɽ�b"O�"�$�AG*j�*�ܥ��m�y�� ެ�X�R7ַ�@��8��p�5�����Ue7aD�&�W�#\F�X'��{|�LW��x�s�.����A�ڨ�#\�i���N�MIi��e��������iۅv��xz
�����f���(�Ʈ�:�X�ዓ��u� ��
M������*6�Y�"S[Is�|
<�������p ��:FkVXf]�[x�8f�H8EC+\��)k�Xq�B_NKQ�S�"�W2�$W�������&w�U������|�᛬dXG��A|U6bJZc|�=V=5�(�W������Ax�k�"�ek���e�t!��d�O=��["�r�&Z��~��"5�#�Ōn�ä���������q<<dW��C��њg�A<A$�]G�E�r��1H��8�%��&[�w�S`<N8b��v	k�̦�ė���J��b?���err�=��>9=�:t(>ř�u�p}�
��hW��}��-�i�P&�n�N�-ةV�b��t�0��1@ٔ.+A��3OQ����5��k�����PMU~q���?Aq$�@���2.��w��To�O��8��S����U7�/�� L~'�ͼ��,�Kw��pA�!�=��puy%p��sTW^�����B�D���d9�J[��Ov�(��]��+�F��W��ˎ
��S&sé�5H�Xe�(�|�a��ώ8�j�jj�L;��%K-pgQd�T �g'�� �a3��8����C�J=�#*^b���豀?�k�ނ]5r��x-�y���dC�O"��L�^�O꺬��[����e+���P���<]�?)F���^�$���@�3)_fڼ�-�uj1�莅]m)�g��9%;GYg,�4#�:�����Z)�gD�`��r�+�	���NpZ_���������T��ʎ9Dj�x�_�"�Z�k��6%3����׎-����2M~���6���_g��Pƿ�B/�-�y B��?}��|� �ڟ�� ���q�䖙�����mt�7�˖���>�nC�͊��ׇg��q{��ݿ�a�
_���nS�N��V6v�'Y.�%��P�ԃ�F�ݴ�a�R�Of���ߏ�m4\���"0�]��55��̱�9��H?_%�4�u6mg�M�������s���b$�г$
�Ul���)����R�B���� �K!h)�x������R�J�� I��9-2���s՘ȶ�D]�a�:j�m���֔q�\�*�jS�.5�o>�U@N]j$q��	����#������t�I�եP�wR ��R̌�.���-�6;Н�ٜ�b�d�u����2$�y�i�钸X���HN@�����0&�����������N�LU��-)U��]|<1V�s��P��Yk�W�oK�cY}��ժY��iEc�Ax����-��
c}���� R����Gms�X�=-\NP�a�,9�|g.�t��V�{>�X��!�rˍ�d�l�����g2�J�앤|����1��sR��7	�X��`�<A�L=����O~/�D^� �"׷]hġ=w.����P|2���D�3��a�/ڛ�_j�M�a�I
��dP��^C�_���Wr����ù��9{�O%|LX�k�f��i}+��K���2�F�� �Ĭ.��� �p�L��z�M��.�?f�T�Fn�j�����f�T�=��p�=��l>�� rF[���_�4d��-G �9�)��EJ�0�ʯ�׾OR�d��'�{�;8>�3e}#��6�Z��=����ç�J�& �.঑㩐�r=;��3��H�5A�2{�w^�(���drP�8�`3'���V�����|*�q�`? |�3��ttz��I �=p�N����F�Ne��j,��Ấ�w�	��{�0�ѾQ7i�qB���\��!�`�Y��z�.���mK�l�(���:�ͪMI��?�$R��(3u��4�7!!5�ؚd�����+��l�pߴn�@��!��2Z�%��-断�	���x{@�CvM7�cª��&�������&�<ɀ �� �I���5+ �7I�������	���>�E�����
Mw�����zz�	�g����_���f�S�cȴ��W!�glj��k!�q��OS94.�����+����t��|6~.��	CQ�Z�iƫ��1s\f,G�vWW��MfbBʼb�Gr1a/S�E��� �v�WP"���}����jz=��>5#ȣ/߉<ѫ�ZH�'G-�ʛD�E�
훡�࣌c�v�ԓ
 �$��,�$ ����SV3�/�-x�1� �++�!1I�yJy!�h<Lͪ�U��7���xCv�E��(���;�'u���ö�C��$��%�R_֊FR(�p՛m��5�5h�i��˺��@��S�|x�iU�ydV�找�ԝ�;��3�"�����J�QkV�<��._����精p, ��oң�H(�� _���F}�83����
�-4TC�I��}��q���P�{�S|og�!���8�6-��f0{$yG6�YRg��I<�l�՝�U�	Q��ś�������k|:tF�GXV�2s����)��i�	 �Y2ި�@%-'O���p���m�96V���U _������B��	su�^�?�w��z���
>���P�/�Hd��Q�-ujH����]wE���Mז���VJ�I�+<H��]��k���Ps�m�a�}�d�P���K�����قo, 8;$��z_-��׮D����h;�
־��~��#��Z�v�\���j��6�;�A����A2`��lSH�7	^y�U��x��o(�b��v���S�^kX�����;24�b�hÌ�uN
��ƌ���Q��ƦR�?6�\vMқoBY�+����y�v�-�;p�Ab���i��Z��2<SR�#'���3R-���߄��L��.�]�5n��אL��,,�-,p��)�,"�%��N�}���젆��9�bCU�H�^D	Xx��	w���$x5ֈ����o�A�Z���$F��Bα���# 7H4�LtfQ�_h�˱D_~!#���Xf��U�q~V��5�D��El{)�9����e4�Ypkp�����7���J|�ʢ�u���.�E����^�W�"v�N�&�ޜ��:7�t��M]f�yl��^�f#D��������Ʃl��cw���jK��1�ߞݼ@gp	y}�O���f��(J��脦���9gp�tj�n�6M�
�nɃ�kK*Q�4ePlb`��9㡥�|���J]�T!�G�jԡ��*ѣ�>м(����<�n�
#�r{��g������A���J�hR�y՟�O�S���ra�3�[�Ȃ�����Y�<�D��څ�x�ܺ����F���+���Z��K�kp�������*	�� �L���k{*=�>�($��Y�I��g����-�]3�6G����E�ּ6`xz���|]d+�%���+B��U�_�6=�����|1�U��_6�-l�r˗���B4R��4�Im�i������y %A�B��s<u��2��Z<*�C�ʿ_�JNL���i��a�B(6;�z�Դ�
`��~��m�@tsKw�a?���7S1s�$�K��[l'���z�����S�������p���dĳ�LMPk��@��φ)qr��	2�UE�; !eщ?��a�Q�ge����r%f'��� 9fJ�U��f�u�U-{�(���6/#�,��M�|��kqy�̜����PQA�a��Tg�ڡ�.�J��t����%_y'����t��	�K�Z��!�MA	��	��r�^va��q>\0,��K��J]�ɒp�W2pq�ꈲ���W���
wǼb��GDi`N�d\�aN{�:�C� a��:Н��@������p�d������K/8*ˠ��Uq��y����y��=���9��D��σ̐j.��`����"�D*�� ���]/�`��{��0Ҍ�(�E�]��8��`��+X<�d���)O}g��#�v1�	E�E��,=�����JM>��Pg���5�}k��[\�3Va���/߮�55���z�n4�p����i�s�?n"��n����4��J�xf�k��k�_.]����į�B��)���@�J����JXG%�c��B�13X�.�6��a&�7} -2W��\��U�3HZ���7��SW?�n�-�}N��Їp�����Q�˩j]������Ʌ��r��s��9��'���(H�0^���:�\\�����|q$��a�l��;b1�|5ӜK�����R����Y��ʱA��֭` l~�z��4�1��-a�/�a5Q�V�b�U�C.!�w�^�̜����qǌ2N�yc��]kO����~������/�{���1(���C�AC��T��&_޹@������o�idA�/���|��!8K�tQ���e�+�20ZlSj5��]�YM��J�5��U2��O�脃��t���y�H˲�T��C�SϑƳc8�{��Y��{�W��g	�+�FM�eW:��Vg~U$TT
r�\J�`X\��P%�����ϟ�[��`O��n٠H�'�&E�jJ�qc��rS�'0G1�%�QZ��j�x�EC!u�z�_[ñ*MQ%�ÃeĬ"���h�� PF�`'	�V���r�n:���rA���<��ٞ����)×w��c�F��6w3�������,_�J��¤��+4,Ԑ����.XO�>���
�U���3x�p7i?6v�fdP��x�xl\�S�D�'}�U�Ι.105U�'�j�B��D���~$M�$.S�x���c����jz��3��A�Qd�)����C��2�FD�K#�@�E���C�V�6~n����CB��	s�P��'���v���w�u�,�U�I7Uɜ�;<l���"���Q�7O�Ʊ�F�3V�>�,ި�(�~>�>)�Xw��C�_��7��d�S�!t��� �#e�0Zw�
�]�<`(]W�"Q&Uz��"��E����V���$���@$4.� �Vy'�R��% �Xk�~�>�GU0�FO�D���L�Y$��LA<�,j��Ƃ�])��ãMMxh�D��Jt9��<;�G�Ug�?ņ�:����ƌ�*�� I�޶m�a�F�﹂�!�wb'A�or�s��(�����`����hN`����谛C~�����ؤZ+�I�"�8����O�ߤ�#ra����6$ۗ��rY�}����Ѻ����¦X~�ҙ�����e�,'4ےI�<��/�h�����Y�m7��I/��#�h#���K?I�:����}g�s�ٌ��G��4�׳�)�xF���8Fw��`wE�׵FyeKw�g���l��x���8�"ha7�� ��6��T���l��4��h�ht5�X���T�(ا����;�[��%�Y���^��%ØUSh�K��/�4��sb-�`@ƀy�)�]�h`�=qz7�u�'���2p�/�xim��7��~M00���kU�baw��
�1P7o�(ou}΃u�܉�v�0�Ӳ-͕ޘ+dZ]�H*��B�\n_[��U:[��Aw�y������ݱK���j�$!"���;n���Y+���x<��h7�j�n�*��ףWB,+���_����:r[ ���,���e��&4O����\��p+��`��go��Z�S�Ă�`���j��i����������=���G�5<��8'u�_hƂ$\��j�:ܒ'��G�I���x
�A�g�#��}�}��V��g�@�qw(]�q8���N����zu�[X��ƻ���H1ev�4���\�eR*��������$x佪��������oC1������	\�̙>n.��G�X�li����؀��_7�=�~i���/P�/1��@.��<�c@�����_R�ts��T=��;�<je�'?Lqqkp����Brv۸��1|�ӶC�$�����1ve�K��pa.�� �t��a$?B4�f0��Ŵz�������;tn		�.����O�L~�֖��C5�����R6��8t�|�t��S�������9���
�r@�ſ:I)�����SM���	�d�~|L���+E,�׀s�g��4��_�Pp^��Z��+�t����O���OӐ���M�{��ar�q�!�`�n�2��JmS���`^�'��f\���'�2{��c���H�KB��\����h5m�5�I�b
��h� �F�ҵ�T{�X�����^E1����E{~���ǟq���|B�ݜ�ܼO�t<�=N�"�GIC� ԭ��v'��}6L�\���vQs�#SA�X9����"(�~J�$O��C��B��/���{u	���?HM�]�������e4�Ѳ+̎�NEafȐ榉�d�:��7b��G%��M�Z]F����>ѪgF"خ�;������^��+q��҇�}���m&�e�x٥bĚeLc��������oD�U����&��db�E�Kݛ��=گjզ�B�ҁ�W�-d�k���$�VqA�`�F�*jiC�eE�El<��o��J��3N�@Eg)�1�1�����r�UcR%ְ8���A�-�ѧCO��Tň̉Ɏ^�<�z_����,1HD��j��U"����;~|�W<_t�V<6I)�����|�,�7��qg�WUG�|��,Ȯ�h��4~J4���w���@ھ
�����n�5S�� ���pHwtft�ϧ�BmBN�+
����'�r���!cG�oQL��䙏�%U��i���v[í�s�I������@3
�H�Xw�����϶.@y�=F�M������)�$W�i���Y���6ڑ��}�9�5��r��6\��pd*�u3Ծڒ�E���U�� >l{�?�<��@��S��uh�ʎ�;�~�XcK�R��Mʯ���Ypjf�|��c9F��j�����^a�"�Լ�ݡ�O>7W\���l3S��}k��<;��zu�;������MBV��/��+=;��`xSBȂo�J)w�.���v���0^.�Igy���|��il ��tcݢ%Z���7T
�R���6�����k���2�r20�<@��g]�ߛnp��?���eBg�Vs[q��L�^��/�جy.��w��JW�,7w1G&�Mb�O�Y;oB�K��N�����L������O�i��A/`��j�0��:�{=��w��A;i�b��΅����ˮ0ء9fj���J�Vk}C���omW��j�Oˁ��jp\L`�U�T��u�6>��v3�z �t���Sj7�霷�6�il�g�dQS�(�F�g>Zf�����{�pl���A��wm��_�R3�@b�!@W;&�)H�pm4�0d��:���N�9��a���͂�_��#�۪?jZ5LG�׬=�ͬ'rL��e�G�r�9�؊��1W�[oZ�`E�s[묜)?��Qc�*1�帘9���q�IAr�NMf�"U#ry: 3��a�JGQ�rb�-6A>]�z��Ac�)�297t�|��޸�&;�ف'R�IP�b~$p��m�`�3J���"P�?,(���V7���"3ӗ|��Z�JK4@���>��ȹֳ�`�gB��!i���$O��e�3��H)*C-ߛ[��Q��W�w&y^X�*��<���'�����OJ1x[or� ���?�P��U��[e��fWﰁ6��&��1�AA;揯'��g�ZǷh��
��[����낋@�y0 �����t6�6`\�l�%�sڡ��BC�_1�E�q�-�<���62c��B7,\�q�ɼs�Nm�^�φ�R��Z��N%qv�S�Wamm��_�$�}�5Y{�
��᎜�8���4:����&���LﺣCˮQ�bӮ�9ѡ�|�n�X˕WU:�d��Fd�`�a$%⦂ڪL�8��fm�$�,�>�� \�v5B�ڒ ����i���Ә�u |	�b;(�"�$wY����8�<z|7�B*���'���n�%Z+�+�x���F��$�Eᦶ%��-�!��B_t�2��ȑ�;�9m����B��ǌ�U�ЖUԯ�Zz�N�zU���P�tQy@#���i !|�f��O�Sf�_W7)�g�®�a�L6{+����� �w�n��nY~P��i��RT��
?KH���{�z�7I޼\�(	����w �IV2�Q�c��/XJ"����M����hX��ĝ��WKL�?޸}�K�e&���t�)hk�ʞи>b�Y��)M�x���%q���0��(�r�6�����aMX��:Ոڝ���dv`<cv�����n�z�s��y.��5ߛYGI��+5Ԛ7���j��5t�s������j}K�<��\x����X�<��*=��a.�ZL�~۱R����b	{�9�r9�C���"�Qt�.�
I��3�l�ҽv?*̈ae�6X0 ���t=��s0�=���kV�b�.Q3�jI�E�`h�Q�}\V`��@��"{��OX�JD<�v~4��T�3H/�̓_c2}׾�ϲT+��y�w�F�RS�{����/`�p��w��a�d1�mr$�D����r����̖�:g,׃Bd�����W%��1@�Ѐ��O�-��r���ol(%9�E�Wl���t+����SVBXހ�=��|�׀2��e��a�o"�^�_3�WYn�/��P�/c�Ƌ·i3�k�f:� ��!Ҥ���Wi�a��|=���[F����xk;�'e�;�S'D���φ�!��!�� �^�դK)�g?_��''�U�e����<���ϫ��PL�V��P����0.�C4uN;>`�Y��&_Q�B�HXkT��H�p���-c�I���>�Ky,ل2��}�H��#�P杦 \��<=�n�$?�Oe��i��"�}�6��/'�2�Ƭ �f�ԁ{�fy�'4A�2��2"�G���K��.��g�q;��w��*�ʸ=��{�)`�y���/�P��%"�.��P�uL�{��v�
n�[lJ�	h<O�0I����73b�F�s����_X+�ڗ�m����*�C���z��s�ovP�_-f�f�R9��Z�@tU[�:�eK�M�34h���~!���xhjN�5kPȮve�{Ȗ�f�S#A����"����O��{����5��θG�W���v��0b>������nDe��3׭�SnI�;��|o�/��GY&0J��NZR�S�/C����+�MU�N��Z��+P-1��£��Mn�_;+x����zq����ȕw��v���q��P�k>?��&[淋�� �8��0m�y���kC3@v%1�OTS�.�ɢ�_��Q��yC#;I��ۻ��ޅY�f�IJ�_�$'K�^�*{/�Qb(�1������g�H��^$���^�;Q-:ߗWS�~���"�S�Sa{�ו8Fz��ݼП�x�5����-�H·����h�H��Kv�	����򯡳}}�d�йI�|���*����q4Ѝ���p/'ps8e�tzB�k��T.�'�TA_t�?5�C�Y^��� �$ �  ʝ��?c���1��ZN�PA��P�3�&fg�9ߌ�W����F�%��0fC��3&#� ��^E%pB��pSA��I�ys�D�Y�
���p\)��a!r!j�.P��P��.�k(H�V�S�*F���]�@�|�6q�ٺ�NU��ʗ���â��#J��b�`W�%d�ݓ���5q����S[�B�EF�7�_ׂ�+����e�+�Ү����V����[���V���$�|c*���?�29�u��Il��;�.���ө�T�:�
��D��5�L\�2פ;�zǡ�c��؟����Z��K��pr�3lBT@��C陸�J�_ؘ�q`<`bp�?i�ٷ;$�`�*u>C�V�Qy��ߪ%��P�=�Atɣ�p�]���O���;tեmb�/$�2քr6F�8E� ���JX�h�88�
O3,*�_}���D����i���\q�>�����;�V�(D���+�D�i�h�X��
� u���T'!�a9���]�<��(�P�ڱ
�q�8�lEO�>�h�Ru���i��E���.�[Lo����6�8��w�N�����erH�m��4&�{�e��~��a�b6f��ȱ����َ��^�'ҋEȒ7L��|�S.�2v?�摙/ 0�T7ء�{/���W�ߜc�`�j�M���Fz��	�[���Ze���t��	\�~�J:���҅0�]b`c���5�IZX��o��~:��Uȸ)Ű&����a!(� V7�~���,�?�7'��)a�\��[qBb��&��`1��N]��7�g.���<Y��EF�Qd���;M�)�ŋ(�u,4�G�X@-��\Eˍ���s�8M�P��t>e����M@X��g	��y�1\T��aV{4��i_�kG	��������d�`���'1�Lq�z�{}�m��4��s����+�ۯ%]��t���&a���懌pJk�9���p��nZډ�<�E��K�V�P��'�mik�k��2��V]L]��BE8Hh�
�SV�O�ș�t	%Q�{g��W~���ݥ�:F�9&�iT��� ��2�M�1����22�F�*\��Jpf֬�T���#�5���0��!z J$�8�h�e9��u�9���^��,�( KX�_����*8�b�B� y9������T�Y�k!�J�j��tG��䙵�b�C��<��]����\�vQU��{���(M�:����'<6��&5c���- �Q*�������˒Q�c�	t�Z�e��v�e��A�[<#dt����e������;����:6�nu�I; �/�B��؞d�
�z�CUS���e��6j��dHo�����1O��t����h�3K-�U1��C�7p!i�r[YX�8,%����c�S�9�E�6�p	�T@s���L�E{���^�Q�l�UՌ[����q#��HE�!ԥ�b%"?i
�(������.o�ˇI�}˪[�=���
�E�B�媃aM� �Ȣ �PY r�WJ�*I~xЃ�3L�J|���C�T	�j=Cz��s��]�M`/y�e��&@L��.]O_6��΁�Z�ݸ�H�d�s�PF,�v#[F3,�H�~Z3�8�ov*��/s(�`m�D���a�M!ȅ�I����4,�^�7f�/�����I��UǓ�q������"�=�qJ�,q��<��
���*@���^񰴲U�A0mR��jiV�N�ncq�E��顎'��ϣ/O�|�*�kmd�bdd��#ч���
���61��n@��߭e�ls�z��80��QD'�4B|7ǩQcg�����jɏcrW]��:�r�(�斸@*��u�H�;�é�ׁ�Y��z��9�1�����x�2$g�x��w���#���p�r�[.f�Ӌ�o�	����-�gz�6󕿚��������sg�Y���cg_�?�zd�
��/��d�z&�X��Ε�Ջ�����C٫8��C@���9M\����Gְ�	��k8Ҋ���B"�m�8�>��pQ�� ����t;ڎ��xQW� X�L�p▹ssc
���@�]��e%!��,b��#�tq��K�f�p�r_�1�7�I���=b��
��rA2I`P>��Aۗ��	����5���|�V�:LniP�Y��#7�r�RD�y��n��J^֚V7�.�֭��w4��,�H�֘�g2]ߙp_{���K��>�����
Y6�����C�e�΄
��(#"7Fʧ��'̵�O��S�֢L�g�k10��4�3�ٮo��"��`T,z?<��E0�Z�QVT�3��wc���)w������K,�,ޗ�#��@�^�q~d{�/���n��hI��*��Flҗ���'+)�sy���	>V�z�?5���t,��?,u��|�(zu&��T���$:'�͝��O;}��T �볢;��e�����J7�,+E�����r����:�ě>�,�a���V�V|�A��s��ܨ�����&�����,(
�]/(,Z�;,k[���=��^��/��cԛ�Q�t?��X������CL9p'��I8��:NӮ!�K<�?R��`�c%qd+p�Nu�S�*��f�&Ʈ9��U�a��l�;�s.ɧ���0/�xo�淕�GP�w��4Qh�{��7�7$u�L��%�(�� ��rsf�{�t�÷Е*/���'��Z��!�Z�0�>�2��䪙�7�wqY$DZa`2�Z�3����/a�P�7�	a=�г��g��(���F�{O<+�.c�C^�D��!�? �/-�o E�O�:�y�#n�i�D�mMV��E=iAH`
ʋ���يY�l}(TD٬���>!Ω|��	�A3{�Bmc���M�PŎr鳀o�4�3)�?tx
_Y�V/�O��㘥�9�(�rWz��0����Ё��õ���}����e��s�	L��'/�W�`�1�޲���i����$����PWk��u�`��o�	rq�v�@4���
^�#X�Z~9�>�}k�i�3v��f�C�k���=�k)-�z]�H�`ܴh�c̓���O�����-_�j��iu���ݵ��F���_�
�|KL�7\����}�� u:/e�/���$��+O�����(���=B]��kQ�e�'
cu��"��	��UJ=�;���t�f؋���nA���)-���b�s���L��lU�ӗa�ʮ>2��`����<
��y"�����������	�u�"d9���K�e�tB��`}.���U��l�B��.C�y���,+$q���o���b���=|�!�ԯnц	�Ҙ���$m�!�:��\,��!2+�b:�[u�O�T����w2D�8�+��洈�S��'��Ķ��9��r�Tz��/4��p.�"Ay�2�Fg6 ?1+��e�Z(�A�U���6dգ�+���s���'~��2*�fEvF���,p%���IZ�|ֱM�_��"2}I!2��>�=�Hz76�/����q�5S�Ά��-���<�?Y�$��3dA������*V\n�Ѽ�P,2]��\t�^6�]ڴ��W�������e{���Ԋ��(J��Õ���7�1�4=���O��3������oh�,+���h����C����p�Y���S �ʘ���B�ȑ�o�ؑ�4����,�7��s(t�˵���`�?��bV�=�Y����S���`7�V���w��(������݀����\�����{�:륋�u��:"(�I��&�5�Ub��d���.x4�΢@X��L	Ϻ�z��/�3b���W���Br��r%��u9;�nYa"�		LF
��*_u�
C6�C2�.0�`N����b������}x�V��ab|?`�--��9��9YZ�{s�Bs.�cwm~�vs��:Y%̼m�e2�R��V(z�$��U�Ԁ�2v�.�R��r�	���� {�oZJ�g�� ^yU�j�ٓ�ծ1�4�������	D��z�cI.�Ҵu{w��gi�&T&W�T�����,����ʞ�ٟcq�⑁�O<�NA��X���
,����K�P�'���޷���z�0��Ժ�U9���Lrd�3��p�$#>��Z��o�.��h�y%e�
�����o�@�imy���U�	��s��u� �es�f���%.k�<�˙�s� �m;�`0�/�˒5�a���Q�n�AΠ���D�����z�z���w���tR�g����ф!$D�a��d��2�z�3��������y|�2[��w����IO�GD�<��/+U�����l᭐h�K��*ȁ������L��*����[� Y�Y���f����g4�غ:�MPj2%�⑰1���*����ۭp�NsPY���?b���I@�������/���VrOS���Wӓ鼫��I��t�//����u���0�zӷ?�o٥[��	�4�۱<d':C�T�/��A�v����=�H�
����=��ez�Dh�٠Z���P�1"���7�(-� ��������aM|:|7��o�KP�dކ�Q	�O��
7��>s�\/�|𴼋��
OX�z���״�2��8����5�H�.z���+{K�a���(_1��*,�Q�Q�Z#�KD` ��y�t���I�Az��	��a؃���٨�:8�]�� #�%u3`�����5͉����n{UUj��7�s��Ur}/�%�"FE�W��:G0��f�1�q�F\wO�;4_�=�tk҅�xWme���'��f	�w��]A,���"jm������kUEg���J��!�5^�Ꟶv<,?KԊ|$W�RR�Ee4CT����~e��p���w0����N��
}q?7L@T�]q������BZ�#4 |�وq��7~:ԿH'�����ޡ�ӣ����m@<�=~$��?����������·��!p @q�0����jD�孬�;B���MDGO+����%�!��cb2�}[� �mx�i>�K!�8$�_���Ũ�'�"2pҹ����$a#{!��~�M,N��Z�Wu���m�-�gps,���+��AͲ��WO�Ī� ��{̮��R��WJB����е�����Q�>������FeŔ7�
��z ���G�P���i�1n۽7�S6� y��EK�ҡ�&Cٌ:� j��f��Y�������C�!�z���6�j�>U�ӝ�N`Q�F:�d[� �V���	�Oh��f�j	�qC�\��\<�q$`.��,�@K�g�DM����B��FH��&ѣ�.E*��3�(�� ��IΘ�g��Ԩ�O芖IG%�RED��I,n��(帱�[>��M�=��ws��N��K���S�{i�r^`	��<��Y�}���X���S��e�N^�#�Rܫu�/�3���0#r���P�e�Lb��	���C9�f�B�Ԡ$�5|v(NI�}��v+9��n��B*ruA8{�Ց���K�R�}�5�O�IW^��5{q�&X&�bS<��A}]A��O&�O'�d*'_a��vr"<��$�X��͎�Kjk�U2���omZ�m�y/���K0�hw�Ւ�B�$���؅GQ�N�h�5aʍ��m��
䨫Å��wy����'26��L�'8�]mk:Y�?q��⾫�g�V� �,�Z���*�U���k�ĥ��B^���K��� ����mM��!���>2�fzU��Nr�J*��<����
w��A�N~�T��������oa��Dߙ�� �d:.\��t�t�V��r��L��j�M��%ޟsWh�zo������ԡt�$�[<C[��өp���hd����L�����[�;���b��9j�>BGJ��rMϦ�\�|�����"c?a��^�}�s�"!�-�c)f�:ㅎ#������.2Ay&�K�c.�+��;�`x���,�	.`lix$F�}��BWaR��tׅ�+��4k��@�b�������w]�K�7unD��iY����VP��詫�6�f77��� ��o��|����������������g1{J�F��O��S�G�]0E�%2Wl��Ĵz�vr�\9˷�uΖc��W���J�B��]�I#�O�݁���u��l����nb��2���x\CU������n��L���<t��8n�+Li0�]x�g��b�C��f�z<V,�ƍ<��' עJBgyU�6�mJ3\�RFݺx�t��z�%d��U���UP��G�f�/�M���,bK�D�^_�D#pj�<��G���R䄔��ƩX�f7�%��1��U���zE��J�YW�>+��tP�	�ْ�6E�)dMu-EG,9۾�A.����I�J�[8Q�|GD�oj#���&C���'�sӺ�ͼ?9�AԺ�jPv���]���h5I��i4���0qa����{�y50���+{�(��B��tu=qڃ��G�@��+���}�bn��_H��w(�q���W�0�0g8�6��;���RH �G�]A&�[T ęViD����J�`+�oq.d�� ~C@�|Ur�ʖ��"�1�u8�껀��7�����O�<�@��^��@�6�E���L6!�׆�qoU���ն�����c0)���/����Ѝ��>�0E�L;��X��3Nﻳ��� �W�T��V�l���	V�Ƒ�g����v�N +�ő� �P���	���nHk�� �$�W@�*�
NlB������f���vF��EK�P~�1��L�����RY@%�3m�|����?Ͷ�x�pl:��=	Ē�"�3R�P�&/.Fy1\\�m�֡�iy�*Y���o�ͯ��	��;j�D�9c2�>;�=V՝�êB�mC�[����`*�+䤗�+�{爺	���q�rQ�$�=qN�M��^΄����aJ#)1<��E�)D�w����[�Yτ���p��@����?J�Q�0Ն~�q �����>4x�+��)&��W�Y6���:�2��&WP��)8�p��6�6$��#O
�H��:���>K�b�n2�������3g����,Iǫ��L#P�^f��O��L�B
�m3�ܹQ�z�R��6T��Q�4�̾� ǔ�������D"iU1Of+r
�c�`y��0¤�7���ߔw�b[!J��dr$��Gce�c$+k�9KhŤ����2��UƋ�+�t���b�ߦs�櫅�NV��M����1��aqh�q��/���f���ȴ�Cή�����+�̟�>��X��9�{�E+�O�.se���o2���6�S�e�ܓ_���D��������$� ��tc�L�é�q��<��,�SB~�T�qȁ��[�C�qhd��1:"�كr�Py\_�s��S�QV��P^"����m�k*1�9�w�᪩�b����IH� �0�K�2uy�"C���P�Cx����nPf����۸_xͭ�=�D�jՏ��P�7 ?e2ݻp�/K|_�SX�e���ḋ]>��r��;e��u�x��������+����S��O����� ��T//�[� ���z���Ug��|��/1�)yiC�)�<|�L'w�V�O�<�`\�:�iQ���BNJ�ȟ��l�T�{�bR�;�������� S���B$Z��GO����H�W.�rXV;��џ���)��_�x��V�N�Ɯ+�{�CTi��:��w���m�W�s�%�"�B�Dy���II��^�U�O�r����r���3�c����%,�
��ﱋ�5��v���y���?�O�}�$5E��׵��X�\��{�XQ
�r�&P!�����F*�͒���=����U1������_�-l�̸���,�S}�R5�g�p{Pn6%UR�x-��Q����7؇��j�?���ɨѝ:f�Od`�S���}��!U�PD{���t�EV��T�h"
�B����Q��OhW�[��?���6V��P��l{LGN�Iab�T�v��r�Ja�d���s
��ӚgPƍ�¹N֨4I
��H\�M���R�և�h�T5�r�F7|�ȿQ�?p�ee�1J�pn���hS�d�����CS����˳5�h���;��q���4��=lrm�r{�}r:z�����b��s���05��Zk^�y�^i/y�H�%�1��~@���Wʃ�WC�*YpYԒ���^�p=�5O��wN'ɐ����{��=�ni·@��|D!��=�N�N!���9gb�b��K�3�-��ʪ .��fKE	[BF��=)��ǈ�!u����~.�eW,>��%�����a����pE�ö��&�t@� a59�`���[�^��ܣ��@l�r@uN?�ƩA�D�x��ʏoɢmVc��B��s׬ i/�:7"@�l�d�K�	�NW@�>K���f5��h��|���1$%�c�Cx���0��/��E&�2�W�(�Ghb�:`��c���4��k(W�)�|X4 `Ba[nߪ�����~C�e8���������A �5cR��h�?S%�5B����d+�e��q������!a�9�x�4�����"v&�P�XH�8�ǂ�l+��|��#:Y=���ҏ�h���O_��[�?:�H�%9�tT��Rc1�U�2��p�.+��p�Yt�	�N5� ?sOe�A��Je��U�҆�4)��@�Ό6V2��]�q�ĭ�h���+�h��R���OUk��n��Gh�1��];�]�}x�M�K�)]zf�)���"��L#�h��'cdw��F�+����m,Hf�FkI0�q���ؔ�e������ft��}'�Y�e����Y��д�&�6f��T�����W�G���l��I-V�OA��x��{�E�����*���k��Wm�ٌ�̉xQ�5�#����S�B%�S����Ac�����>Pl�o�iiϢ�T��
͛s��)�_d��@u����ʩ��bT�"m�X�Z�[�B'B�>��aӋ.����`S�#Q2p}|:�N xjFɦUw#��a�z��LZ�Y*�Y��p�50?�9U�$���!��+	��h��?8Z��q�$*�Øͦ���w�9e-�W��^��+��)���z�;��5MJW�����"\QBsAoi�����P�r�яcu$ ��Kk�a�ߩ�.���)�܈�#A�I����س��D�@8�9�����Z��-����`8�~d?��U������؉W)�-/%Y����H/7ጰ暨	��JH��8��w�MW� �J�5Rbѫ�iG���tQR̢�"�C�ʱ༕4�c����{R�b 0��S3r����؅2g��u���i"�tN����mJ��kI=\p��	ӽ45{q����rL-n�$|y:n�U�4��&�$�I�toz����oc��S*����PTU��AU����ey�c��,b�o��M8�вZ�Rx�jd��g�Ge#�q���ʻ���sf8�3��}w����(r��}(8�:�5���ө6Pܿ^ʻь��E������e�~���¿�F��y�ԣ:���c�rgt��bY�%���b��!�[�̅6���rg.k�a�4����f�9S��2 	b���ޘsٛ�d@��NM�ҨP�e�QIF��y���OCV����;����$;5�V�����	_#��MhsD��7_n1;�38���	�%���g��?��ٻK���i�{�[]�u�Q>kT�r�P!/�t��2e28�1��]��&h�xV{��8*�b2��P��A>
ٺ�m���/��n�{�MK��]�"2��	l8�P�|m� ���ۯ�[p�6�6�r�1�c"�6�viU�OI�b�oM�fF�Z|�t�F���A����^���˺B�e��+,@L��槅A������6c{����/�|��<�Yv.Ǖ����/�~٤X�u;��G}E8�B������pL�Z.�=5T�giV.x�m(7���-,�ס\	��P��b��̈́l��p�_m�/t�����~�Y��@i���r��W�A<�"�q ���@�N�+�����Z$'|e�f�t��x	�f�Eݯ�B�s�c]l��m�)�,)rׇ��sqF]Ó�a����DK��[��.C��-Q���f4�F��
�����/z[�5^pC<�om0�vyJqZ	�f�p:�i�e
�"~!�p��O%���e��@:���@x�Vm�����`�lC�c�,*Y�t9b0$E��v�@$�[�~��`g
)�i{�+����r%�C����H��q�_J���o�,@��G]�|�Poi�t\��"3���%�j�D�{ ��k�	d$>s���?UG��j�vѳ�c�:.¿5��OϋU�m�8��lUص6�\��:�����DX��E�}zY��C~/\L��
J8[�"=�δ��j@���0��đ�M��r݇)M����y�x:ojl\��'���������.��N@�Ԙǩ�{���Qs�t�\�jJ��
Z�L�g�x*3m��M��$ֺ��e,f�W[��2H=�:07�ǆ��9I�݃\�ή�%o�lN}hZq�Ķ�к�����C4��4 �#�W�i�]>#-�:��V��-Q^�5�L[�.0~�Vu�d�h��VW!i���|S
x��xX>V[Ԇ��
i���6��o��))�Ot%��J@LyY:x�R�}�̶D�m�����"��?VH��,3f�xZ��B`&��q��O�bձ���&��L�sDi�}!5��\�0ҷm�@���n�S�F��b�oe�V��x�0�% k�\��:4ݾ'SS5Nդ�;7���]�
�i���x�oI��W�^�L��ŋ�"�� �����|M6L�PW| 玌��?:CJx��)rD���[~W�``������bOQЍ��,�6w�u����MĨ���.&9\����?}p�����5ͨ��O��#Oj�nO�wf�p}Lq1��X�ݎ�a��5f����4�ψ�
_#�.w��	9L�dO#��q�7ڗo��Һ�h�un��ۖ�z%��g�T�Ή,x"E
'yݢ��v��r���1���{t��[��ׄn@�c���\���X���֘�*\>�㑢0t��B��A��("��/GcK�X���+:3t)sJ�:���	+������#M�J� vd+8v��!!��S>�Mw��}O>��
m��z�\�%���=�� E#�^�"� Խ�q�4��Ny�)�4�F�����+8j�vz�da�O���X�;V��q���t��>]�A�>�a߷'�/&���V3@.4�&&��� ��%�x���&F;Qx��mME۱�]��uݩQ-S"��10�ɭOJ>��":jX��R"v ��y��ԋPF�й�DZ-��wp�����&p-����h[�d��t�{4�R�����2��yJ�f�b[�����	���!�K��,S��]�Y�3��p_)���G��Ү�5D	�5�Lqu�T��n]��C���)_&8�~�}r�(�
��3��I��Q�ہ6	x�9[wp���>MENK�G�/�{9��,��>��!n\�^$�_k:'+U�Ǘ�����mi�key�C�F�p�*Q�f��h�~����kDS6�yn��hs�:0��j��-��
��f�y���@�Bs۞bvڴ�8ئ�J��� �9񦡅�Db��}y��%:��|�)��y"v��pA��y�6Лx�޻� "_�� L��㮠������!����YB���k�㢊v���ݦNq-@�
+?b^���Cp�mU��J�r<�S�q$ۑ2��-�cS�|�Y�NB�y斌y��r�u��������d��ƒ�x8��#�͖�T6�v�d��c	�	s����j/������՚�V�wb9��ֻ��(�ޱ0�%*��	y�I'7�k�LW��lL�#�~t�N�-�1;E�T�N/�I
Gk�VͰ�n�{R=jo����yu�
����d��~w*���b����}j	����e W1v'Z����.�	�<��,��$׼ĝX|L� M��M�E�}� ��lq���g�+�䴖����Xp���{!��͏ɏ���vȫ�g��`��1(�q��X�P%���yn��'�����M�Кh�׈���m���_�@�����J��ŭ�k#9C�B���Ѵ٠�Zt�C������Q�#�B�տ��C�Q_�G%�1�.[���V�~Fm�$���aB{3�l������^�i|��tО�Kn����u�a��/W߹����'<ְ*T%D�m��Q�.�5h��B�����*����0�9ry���Y�E{'��''��f�V)R#�5�G�	�T"�[�x�T{��2ܿ�X�Ԋ��ss��??K���#З��2��R�*i����a���Ȃ�6ɋ�~��-��G�<��=^Y��$�߷�|�n���R�إh�yM,&���:7'�-ć[���y$zq�D�����!��� ��|,��MuV��A��xB�l/Ҵ�I�7m���c+N��'�%�uP��k���@2�&������(L(?|�3L+�+Os��E�:��
N�*��-.�А��;��Ia�^�����(Wb����b,���n�OE�̐d�'�I!pJ~Ը�z2a2����n�Ip�����}�]��
�5�0;��	qq�M��6e��.�dqg�L���91w�y���p�xs�q̈����=a�]�Nb;�J�5�$Aڱ��r��ҵ��4��pK��(�ԮG]rJtPJ6���[�FTB+�e:��j��0����p�B]�C��q @��;����-�kwce����JIr0"�\v�>�0���nJ��$ÿֳ��p�����g出w�/�vm�+,�}���V��ߩ{� ��ɕ��l���9N��\^t��ڄ��̦}�v�&����h+ma��"�@K� �Ҙ�W�<�����H��t�Ϙ�;��Sm���\�ڼ�~`q��d�0��􅻸.`�(m��m��{Z�s��Bu^��?�'Ч��d]�j��L��%��Jy�>���L�Zu��8�4P�%�8�AA$�r�=|�0� _S�d�UI��#B7�6z�Q���ˠ3w����!�tz����zB[��ZV&���wd��I�j���o�!��q1���KH }6|�l��E�;�cb�L���$N���hȱ����z�ew�x�����io|���'#c�&����6HY�١D�sDat�r�x]։�[1K����Jq_��	�w-%n�ޏ�����x����Z�)��b�]Eau���♔5��n&T<ˁ/U3d�e�W�+���%�2g���wĖ��x��Ɵ�}=�0"c3��2&�U�M/A`'(T�ś�����[���e�Y������rtN�h|ݘݷ*�gc�|����������%����l�1���,�鮭1w��~W��} �C��%�KP���yjMɰTnQ�f5?�|���o@����(��8�Ս�%�F{ �G�oI_�+x^��D*�C��PC>ʧ�b���^b�KQd`� �Zx��w�f��PL��t�l�C��/�8����;��y������8���G
�p8|~,;��ܷ�?���
Ǣ��z9�I`�7�Eu<��8tp(�{D��,�i��D�k����jwM��HfK}3��xY'0��c�����9�h�\B�!A�L��s+��U�J�vq5995��1���H���U5"�Qz��Ou��}��P�N��+W/yh�����uXAz ~z=��@f�7)�߶�'�jF�_E� ⭁�@8ܫ��	=}���e��������ŕ����{�,��? ���|���qVx����N3�Z?'&vt����z��cs׿�Z=ы1��MZ�G�����l^�B��;�����w�\$ٗ�-|ڴ��n56����AQlch�-��"1�i���������~e�d@pO�x""JwRp�e�-��s�����g%N�c׸r������[�����)?m�-0�_as�̹5�������\a�9ՙP����/���< �j��.�a��<�tC�3���� ��nˇ�(ӑY�܀N.N�k~�xUw(<�k��l��d6n��ϛA���<�����1�7u@Q���oU�{o$ƀ�s��޵���5(X�A�|���X���\L,��Q��u��k�ձ]~IXp�8�Г.�\W�FQ���~�pY��>�)!A�V�!�w��$��ԡ�(|��~�-��CF�i�ǂ���uاt�B=���mv�Xg�k��^�%��]�z1��R<�m3蟻��4"��UjCn64�|��[d���������y���?$
ýfsf�"�V��wbT����K�'1?��Ro�y�0i~\{�J�dHF�5IQ<�^0νI�V�h�^�"JK݌Bf` pX��Y�<�H�Z*��
?��b[��B7�����xym#?�fn�}q��ۈ�1��4��:_�?U��!u@�W0a����y
���*��}/:�!{_9w��L9
��W�-XF-k#M?p�D^5.�h���}UJ�X~�oi#C��z��������9����5v�J-����@�Gu�<�Sq<?�������5��x��Et�O�r�����	�xo��~�n�d�~cŎ�L�_9[�wBQJ�=�ְ>��uz!�'ܗ���9p��/a�2�_�9)I;�:�"��D.���e���Y���f,�}[���� �ϡ��	@����"P��(��8e\�wV[;:�m.�D�Z1���{)ا�d��t�٪J���2ˑ�����;Q�'{,N���R��)Z��$>

���dF3��/���d �6�5YV�+Q6[$�z�`�pc�$�pqlgߑO�]y���,z�Ie�]�/����\�f���Ʈ@j3��Q)u��6�P���)\��o��;�9{J=�? �$�7�8������C���N���0�+1���w�lp2U�K³�gw��U�y.l)2��"y���G�^����O�4Ŋi�Y]�Ukh���M^"��q�7Ȍ~��H�$7Ĺ:I�����#Û�d���q�`����DH�C&EKo���ٯ����W<��*&�uJ!���g�ž�D���&sU��X�q�8D�KD�|0("Nt1���+Z�/�E��W�]�Du���+ޯA��XU��%����d*��ȁ��Ր���S��U�����V7>����(�%�����E��&'�&Jj�:W=���w��P���5ʫ���C�{X|��&�*IZ�k7?"�"�r�5�r�>FC���I^O����qM]Դ=���#��\)��O���&q���2�-g,�θ�k���{hד��P���X�r����@�������{��Wv�LV M�7��ľ
v�qz�5|,8�+��P���/�b[x�Z�"�>b��Æ�=)��`����\|�itw��� Ӆp��f��`����\�ݒ@���k�P���e���3u�j
���s���3W�ꤘ ��{z>������W����z�EL����m��󪄄3�M��ȳ0�n��VQ��J����a�G����	HU�h6��Ȯ�Y�@.6׵�ō3vxs��ΒW> ra,��AFxbss�Y�<i����t18�CC)����z2&ʩ��[��P�히kI@O�W�K�MJ�!�k�c��QJ�b`�4$��	^��z���v�F���(GKA*���8_��frl����k�8�:�������ӈ�G?8,m��M	�#�U!޹��{C�x]:&g��X��w+�k�%�(R��,]'�݊��|t�t�{�ܙ�0��u�}��1q�16P�V�m-`�̠�n59@/ �m�u�~�sP�\k@���	�9�&:��4�o�A ������[���E���U���B�㰹"�7L���0��!�x���6�k{c�A���P�w�	7����	�Re7zy>a�_����m���>#l�ص��u[��b�����T����6����`hϚCG�+ N�+H����T,�y���(XJ	>��o�sHe�����݊t���1�G���G_
$u�f!,P��舱� ���a���kc׿к�}n�
u$3�M�T��޴@	X�v��	?��������ω>3��9��^�
�A�U���{��~�#/Z^g8�H��d(k���LKk�W�r8�۩z�X6N���2�RM�<�;6�G����:U�S-kh���)���r��aﱭ��݌��-��u/3�2�T�(�
�ͼ�@y�ێ�@u�P� Z5�r�[B��t�~Skpj���J���oK������<@T��m�pF,4��0������9<��q^�|X�ê�q0�r���a���_\|� ��x2�<��0��	F�<�4�A�W�`�*!֯/�3�%��T���'��;���C��s�ޟ,E�6=���T7�C��������^*���Q!Ov���d
p�I�Zp͇E�œ���E�C{k���	&��V��Y�w��+܇S/ٓ�}�� ����3Ǵ5��w�^�z	e�{�g�d�T��4\�p��B�:���*H�]�q:[�V��.�������'��B@8�ך���M7_�C�*&�a��t����θi�z��S��t*�F=�fTTb���A�Ĕj��#=y�1���Y�v�X� �B�mc���O h�YD��\h{z>+#��BuYz}d ��0v�߬S���_�pBe�cN�ܛ1�p�-]R�r6���d6�jv�Jµ�k������ښ��������ʛ\6�I^�5l���)�+X��R�z�׫���#0�z~E~`��բ脦�d���Ҵ>W@V�?��c��gNW�69F�b�'&t����C�:���I=p��>�F�;H}��x���M~��f*rٓ�f��hV�3��B=j��o�Fuo����	�"
;aZ�����[)���-��4[{O�b��{^ˤ4}��|!x��T%d�1�:1���Ö07�p�%��j������-s����>(b���p8,�&E�n�$�^�07�.sV�t�g/$Q�k,�)��他�yrN�O��"+����?��l���U�fr��]K2� 5+߮�vʆ:�Qd�k�梒a�B^�Ռ7����̘�Cfв$����M�݁����g��)���#i�Xˀ(O�涌'����=5.���G����"�`�E}�Ng������Aؚ��@�،�9��ӹ��d~���=�c��)�m�"��e!ﰹ�q"�Y��6 �ް�@��!j�TJ���!�J�*�ݺ����,�*'�g��rĚ<#�s�u�b��h��6�gZ�_W�~���q1ln=����9� JV�$͢?t��5hU�=(4X�J؜ƨS��m�F�u�(U��(kU1�*��S�?�����3�=G8�y��N�j��Q��=�Ӡu�'�Dy2`1� ������	I��'o� Qi$ $;[f�َ�A=�z��A��o����ܸ�5�o�4�F0u,6�6�04�;���Vx�Z����ϲ�ϲ���SĒ?t0���	��·��^>��?���P����:Y(��Uv���V�F��I1�z���==�����NU�e]ʁ�_��R��CS�FG�w���x�Ѧ��z#�����gM3U[��i��l���m;���
&@b?�E�u���;\�ho��s0Xze `�G����gQDnXl9�B����Ɔ?�[/!J����u��2уふ� �g�.ގJu�o������V����<�����eg�%�
��z��ϺF�%�&(L�7P�;�>L���_����N8���2�y�궆�|I9�"�(�����a�Ư�@�Y��	]5!��%3i;���"X]�K�܇�P�a�wS�*T!Y5�C�se>���vg;�?�.����+:��lt)9JTBS+�>E������Eu�T���i(�f ��=�U?���.���8,O�j�a�
����TR�2Ft�8ŕ����#z�df.[vu���T��۝��9��r�x�׆;��	�H����E��eb���J�>��&��M����)P�/>��|�1�qu�(M���>e��T%�����r"Eg��!4QD�\&D�2@���̜��y�Xk��-eVf<�nu>7���tkc����j�R%�"�&/�)J�I��r������R��!�7�=gcg�/����"|-rR��ՠ����e�x���1�DS����0�����t>`���M�%`����.��ʊ�l 6L#z���k<3�hjQ=:E�}S�jட�+'T'ᅫ��ա��,�������A2w��-����fx1�;�x�l��Qx^pn�C�E�j��+�Q�Y$��ߜH�4O��(;��V >Rә1j���!�Hl�H HaCN��ڠx��S ��k t�;
9F�i�[�0�xu���\��+1m�*b2�� 5V]���R���ӵa��pvN�H�Dr��9��~HY�on�M�_�$x��:��/���}��U~>dl\����Ja���jx'�Ғc��p�J�!p,�&���C�[a�~*X�bDVy�B���WI⪠�j˻���J��
�jK[ ��P�X�1=^������>�R����v�V�ZńӨ�/��z�$G�k`��6��,����|��Ƈ@�Y�m��i�����-3�Vۑ8 �-�{u"�:]O����z�GX�&GT+λ]�XÙ�Ƈ1�.|��U��1�a`�JIq��ˑ�'�\�J�8~h�1{���N��s@��� L�%�R@i�7�wY�:�����29[/��(�����I���f|��aj���@�u��,��!��Wt�'���e��;�\z��ZgX=T�ڂ��m7]�P�r V��5�GOB�e=�6�� <�����m�'B�:�ggsS�ZW@Ʊ�Y�O��E���@��D��@z{ȣ�Q�\ip�_��_�rd4�؈.�x�6P�c%~AX� �im;��^¥��"!�A�����=M�Q�u�GpiX$-*��G*�|���J��n�3cN�`)|e
&�8, ����m#����(ϭ��V��*Q��ʕ]�5���&�Yf��HZ����\���I�����-�TN1��C�F	�`�����^�G\�(�O�i�����G��lto#��c�,��?�8���������ЅP��ڧ��Z�%L�׮c�;v�A8Pｺ(��_�	�5�`�yO��3��>�߳��h��Ŗ�S��L�m�Mc��BH-W9xF�5m��� �Ϊ��:��f���$��5�
S`T�L +]T@u��b��c�de��E��_4޷�P�7B��{Tsz��&�����A��	K卍a��ٌ�k�-i���߳�����u8��=Q�2�����v�R�7�_wa՝6ƧI�pzJ�g��ԓ����UQ�!�_�̟!p*�k����f�kܧ��!�͎d�@�"�Bc��H@��d&�Y;cܸ�|�_�O��wp��$*��M��~�����3��Lh˰h�V��q����[|d�Q@���6az�ˬa��8����ON�$�yMyU�����$P��T���^��)�04 �/V8엿��u�g^��9꫿#���܃�q����8=��]�f�=o�X(}�61�1�O����Ћ��u�6�,��붲}�ۤp��FrN	r�&�]�ۚe�><&���=���*ym����������K��0wY*�4����)P׻\W>��w+����)Xg栈�i� E{�L7'���5v��en��g?�`G��i"�<�S�������������k��n��Q�ɗ:�#2#4�ya�L���?�kA�C��Pַ���]4��_����f��Q��i\�˩���$��92�����׏����
��F���S0�1�y푾A�0D��'�9�#���e\�ZȐ{LW#S�F���=��]_
X+�V�T�Sx^���։\�����������v{�.�g=UE�)ɢ(g��o�PX�_EbG��vWq�p������v�Mfʪ���|q�K`��uJf�ϯD��������n�#�"]��Ǐ��W�B/I��1��m�G��з�f�x�/�Rc��,�˵LUGeJ���������!H���^P7J<�0OS#�+���{/U�{yJͽI������ncga�r����2�v:P)���F��a���$1�HJs�9��@���L�0��R����So�Y�)����o��k�w��#~ ���Yr�oIXhI��hkG�XQn���t;xP�.ZM�jX�|ңI]���i>t�Z�<�8A�g���<?$���@2F�T���_]EDK��������:۹Nx�TV7���t�l��,/!r�Z͡o]���T9�P�CH�wZ	�>�u����д��3�H]������ <@����j(����^��O>�7C�D�J/d=W���R���b��l��7��O���G��)C_0J�V��
o���VdU��A�!��^�nv/��(�j���e������a�� Xh��Q!�ey�_��r���t��z�}���zn�)�� ��vE�ق� �C��B��R�^��]��Z��{b�j�6�)�y1�P:Fi���CB��q+L\�n��Q�h3��6$��.���8&� ���p��@çij�B����G�g�^���3�e]:�w
��ٗ��w~Wd�U��Ԕ `W����^]��(�4��;ר�i.�ONM8!�,��ҭ��(H�%|�|�R0�Ԣ"��r!�zb^@���/W8�_G�|Pҵ����튥�mד>eI� Ժ�{��)b�&1��B��"g��A�͊�ً��4�*��d����c�Ů�	$/�
�����
�(��fS�g�"h����
��c��o�nt|��H:T�q�b�Ό_(��uZ���h4Z@3y�^�'��Go��W��U�k^8+�Jui����o��i"��[�y��m��9.!% �%nU�,���=&҅F��c�x"d�@�����"���^mek+�`)��xT�R�g�ab���?^I�
��n�"ii����V#��+
1nh�>g+{2&c�� |a>�h�M��9��Z�]�y6Y��%+�_j9rj��fDI�g��ԯ��~9�[��)9�A�H-�}�y��q5��<�M��^�BR�8��\��7W��gih��ij���3i�㯫���o��+�G�K��^�;c�#MC�l�G���\)T�	2iK��
�j,�^�L�,�����CD�����L<���>^dx��%�.�2��s-XΊvv��@���^P�bUt:19}�����+��6�CB�v��I;�tx�c��ǚ�,��@jƕ��4�M?fÑ����jy���?���{��1m����O�3.�!C�˨1�!��h��4t}�h����}`Љ�D:�@�כ:���H.I���p��~/ƻ��k���.p���BG'nz��������F�������@�NF{�I"n>|��2�-�d� 5�-.-�5���S�-G�X��V?��jW��켁orQ%������tD�fvG�mRy{����eE��L���Z�8Z���K� n��j����*�`���&��[��w�:U�Fޗ�,��+HB����Ѧ����vd3%���Ah�Y��R	Pi�F�*�◞ll�K�4�߯�%��5ǌ�M؄�q����. �����ɧ�7�ޗs�]>��7c�1�a[w[�G)Zw`A��Ѷk����H2S��V�}d7��h��V�&�Ă��<Z��kD;���۞�!�yal3�F�y	5��H��b/�IZ}��Z���D�Y|�G��HcW���L�IWܫ/T-�	l�7�Ze���b�y>���Ŧ�P�ȇ��Z���Y�-y:	�e���p(x_&���s&����fy2w�L��sr@����W�����G0� n�=�AD�FUwo�<^�%'d4��Č.��Z(t+�T�l\3@� y<��L��	���� ���4�O"e%Z�ܿy2g�|��,��S��.�;x����� �:�L�����%HJvT�����%n!��7|�CL�pzlvS
dCs���S�Q�*����m5Kj���k��ƁzzS��W����[g�du�w�e�9����q�E��5s�+a�D�t�V��K���4�gN�ڱ��W�g�J�5���˶����ED;�i���h�pK#1*��7�Ҝ�Y`���9Cؖ����8J?�7H`���kI8U���j"c��/���˕�ɸt�t/M�<^|���ә��uY[WἛ� j���F��˜�'�i�� �T�$����O���$BH�q*nq�]D�3HaƱL-!��U�_���G�����a�*�7織E�rJ~t��N)-l`v�8�]r�k. �\yȒ��Ƅ������:�G��ezg!1A�|����Ar�d���Ӌ�v�p�������R��LЊ�uI+4�f������T�q��k5[����#.&��3v%Q_S���d��}�m�S����E��R����M2$��6Rl�l�x�&�y�+��C�L����E\�3�;1%L��\�I)����6g�^a��W���--a S硾����G���H�������޹$�M�W՚��]ز��?ߐ��->��h_�a���U!���I�*x���;�;|�]��-�%��+Cbۇ\i���x�5o!o� ����.�MVJ;3��R�i��dp��w%v�*���=���_\l���l���j�|��pݼ���P1���a>:[�����O�U'��Mس^J!!uFع ʲ��R&ݰW�q=�Ƽ���9�J����.C<�x�<Gn�����
e�ȎA7�c�(0�W�y���z*�vM�Th�>��
�yy���Y>�}��s��I��`��7:���\ ��y�A�̿�ހ���4����y�Cm��RO8ﰱ�ܢEEβ4��u�O�����i�Y�Iw���ML���I���*2Px���U� bt%CIJ������=>�r�:�oϷE����+�lr����::�mP�����+@͗�:z20+�z>���<p�\w�&�|����0�����𙶯՚��B�t�,��QĘ�NoR��5S�͢�8�j��2�c@��fk<k�&�ኸ�	JB5'��%T[��	"*&�4H2���),��3�Q�E��+�"�L�ٗ��o`d�G�(��!Ɨ�nԣ��z���CjM�1'|�m$}���Gn�l�؂�p�zסs���VG�t��O�6ҟ��3 !�$3�Y/;�<��β�":	vb��V$>��_��q��R�������H4���?<8�y0
(��rȠV���Ɗ�Os���|�/��U�5i�:BzjEb�<R<�ʹw�&�`��Y7���;��,<��A�H.mJ(Z%�Z�Px�Ke��(G�4j<�c��됔���-�����	u�jD0<�������h���,N�B�銋��j��*�����F��h��Y�`��
l> ���ȳ\�Sx�U2�$x'	��J���
r=��XY��}���@��=�=DB=���}�T��X��P�^^����Y�u�)�cq?�����("�r�K���KB�M�GT���r��sW����	�O���Vf4-��	�B�(IO��dN��Gn��f��`Z9e)�-�I��S�ie(/��a֠tÉ�p��?��lp��J�E��ď ��O�ூ=�E�d8�o%V��	{�TUef�����O� Y�ݖ�ǃZ:���W�Gk����qH���nd��s'��94�fð�����K�q��	+ꦠ�jM,���JW#*�N ͊��o2P*S�m�Izq��\���7!M&f��7>��n���I�c��0�#�~�q������<p7N
w�v4U��Rwm]X�|�2�pM|��m�)�~3�yC���C�I��G0�2���r�o(�eR%��.��J�y]T�0�cQ� ���헑�,-� ��2v	�1a���+<xM����:��	��' ������#>cLR�$��j��g���3 @4�{y��b,P�]�ꡧO��ÆIrϟw����:5��1���4@��Nq�#sI�^m�I ��3\g��FY��I�ި�;�f��	N������Y�����J�y_�'��݆���C�|7�u?�΄�G��
���[�R��K��Pǂlu�+� ��>�4�<���AL��F����T
H�ZGME��5&Ba���Q��JD�Ds�(odt,O:���;��Y_K(���+�P�7�`��E�b��7F��f�m�!<�I#}��x�h�qTIvՈ��CP��Ns��m�u��������㾼-H�a
��%��u����]����G:.m�g ��?�e�H�A�/�?�����v��0L�H��$�"w"q��Vhe���Yl�
����:>gM�o&t����*]�Z�p�Nj�	�j���A��U�TH/�I�5?E�L��\��c�7dc�)`���\Ǝ�Ǽ������t&v2���~�2�"�Dv�a��� �/�z/�0k�2f���/�m[`���Q��~�
/����$��\�a�^s���`y��I�f����M�wz�5�ǂ?������#E��p�>nf�`���bm���m�%�U~�;�S���R�뿞�;| �n���v.�M��\���m!��°�n����l�����wY�%g�>�~��>� 2�_�YQؐo�����Y��Σ�4=F�	xd�"6�1��	-T���;��U�P�p޾����ʽ��� #l�N����^�?�_��Y ��I�S��Q��i_��h�k���_ڸ����[���mL�Q�L�J�!Y-�pXB�.����"1a���	���0������Ζ �$�MX�C���~�\+{��J��ww^�.�(����$s��a2n9sJ/�R� ~�hO��ʟ���&���Ze�L��K�f�!I,��P���_o�p#��_��p�G�J�Ci"B�a���C� ��Yt�3�|�}��D���ֈ��@��\t�����	֖��n
�������K�� ˎ��e��YR��i-Q��w����$X��Qrd�Qt�TK�F�<����5n�MSx13�{b�[��#!L��0����:�>�TZ`�vb�������S'���j���Ri�S|@���k�>�0�ݶS�����T�ٝ`<����[(����FXz+P]s��ݤ-S=�8^�9����g���H��������K�AbQ��x�fS��luͺ��#�)ᶗR�M��`>��[��?�� [UrR�8���
�U��:�xP�6����<���#�GX�"�ڹ_��
����w����0�T71 �ݜ6��K�G��������n=ZQ_	�0�����톋N��HG��W�r�$�<���%"��Cjip�N*��w2æ�!J����]���|� ����u�]�����/"
�H� !�\����ۧ�S���c������A��Y|�n��q�����]A��l{^��`���6%	1��Rv�Yc��l)�\Q���ļ�S��kx8��خD��RP-�r�u�*��>�L�`q,QH�J�{K]�*Y9[��?YU�X��/Ƃ�ǌ��m8s�Ӕ*q2�gA;��V����wdc�A{+i{R{��9�/��V��4��`��|�K.(�˖6��Qr��� �Cio��P:���]m��'z;7�z��huTDp�'.?[S��A���nG ه�)I�e&���T2 �<�	ծT�P��n�`$^�܎��j�2$p�g:�E��?ߟR�NY��vzcB��)�u؂���b5��L}�����Ea/R���#� ̻W>w���D�HD�x�ꠐ#�J�#���)��3��z�
U9�A�TG���a�n�|r�1�|��9Tяx�������*����r�Ni~W9K<K>
L��s��`��ɉsM����[�3�R�
��&,�J����:��D�(���������|i����9��(;���q�!\��o��q�̿��t��(<�@������=?qh�0'�+���qZ�ͫ���+`��Z�%{�B���>\ߏ�f]C:��(�p�n���H?
(ZN�|;���;�g7��|I�o7X�t	T^[��dSX�?!�kj������bP����ōx��)hR;�Bo���ʭ
eW��-�^AQ���J���H,>&�)uqH\7&+�����b:����Dk�#�_�7X�hu~�럲�a�˂�Pw����<�al�k~��	���� ��"���=���0:����#&�x��&�34'n�p e\`
��>md1��L�z����6+���`�0-t �ҚG�et�S�~֚�(�%�1�L��8����X�Vq���B��<xć@���:_A+���(򏕖��O+�������x���N]S=k�C. ��VkY_�^C��0k�S;�@��&���1`x0)tP-K+�L�~R_����SH������%�*�V���QF�Px_��	-[��.B���@A#�Ɯ�d��f12�Oh�rB&��)��[��\�טڴl_��D[d�rDp��QWtVV�>Pu���։i����G�*o�Ά�m��a�jKΒ����z󱖔y�IF�������s[D;s ��W/7kh~~�M<�����U�Pkv[���=0����.�H)��y?wp�,l��T�.I[} Hl
5-���ED
=
QWJ����p�Q?n·!ˇ�>���]1�)� 2q�Z߯��<2�c���z���"?t���I%�p��A�}���9\av��=��#e�ڿX=�b�\G*a6��F��L��GM��H�r'�b�$��$g���y��c4�	sGjV������0l'C�Qd�c�M��261j�Z��Z����u�v?��H�Z{��K#�WԤ"!�sy��N<'�Q�b��q�¯�[2�\�~x�1����7�[��M��Lh���뀦4�����ʰ����w�X'E�q�+��f�G}h����:g���hc��8eyf�wC/ɉ�O��%Q�s.�s�X;坌��oL�<�+���<~�2M��q�v.zi]��{.(*4	''?�?,��~��n�	����R�S:�#�2�ǖ�15>��ja��I�K�+j�F�;��@s�1�=/b'[�D��״Χ�s��/��tWn")���V'����X>��f���r�= ����� ��R^�d���/k0�n��*R��bG����İ��׻M�I�2_[�k��βI�ԬB�-����p���o��&���J�,�z;�w�1�&e_2��ʴ]��Z2�I�!mc�
A�tU`�;L������) W��$5:
B���Օ��kA씢֩ɺ�ح*����>��($�*��D&]����-U�IT~|�����)��V:Ձ�LY�ϿO��`>P$��o����P/Sjb�����ʋ߷_�a�8�����U�m��<����\��c�U����H��4��#Uʿ��1�׋����pb �#_E�&��m��7?n����鱗�:�]�%����_ �%��`��7����:�/��(�`$Ͳ+
>��6�ۤL "g^�pC��!�S��V�x�w�_�?��l���:��U��A�?�`�谾j;���d �Po##�<Dc�U�P":	��Zd_��k�U�p�e���Z��F���D�XR?�!�%��I�y�:+dCB�:8���VC�k���'���Rѷ�	�8iꐲ0��^_v��'���o�Ή�
�`h��xzZv�~W��*�L�
��gi�g��:�k\zg@I6��ᾥ�nXӴ�B䔍��l)h���Դ˳ e�-��͋���3��F��I�j�;�� �A����5�n�=Q����kLJ�g=npDu�@�hx9�p+�o�i�+Ugw,�ܲ�l�x����3��}�ݗ8��O˵xo<�e)'�,��t>{C��#g���B�Z�K�e]��4���,�cA^]gHZ�cّ����)�e{gK�O	E ��U2!JHR޶LN]PRAk��r�hYj��������:���5HS�p1��t3i�X�bЂ� �ꑘ������PEL���*Rs�GT[ƣ�aְC����ܭ�T[��7jv�D�u�(���CF�F��9��#���Y�J�^ⶦ��r�o�*
�T�Q�
 .���6�^p%i�?��Z@3jj�V��H������3`����Lvr�!�v��7��}~ǳT�O:�����j�5�D),M��3d%A��i����rS}��Ւ����2�	QP�I6����ۨ�KX�v3���}�۠�-O�ǘU�%,����K��x�Ak�{������\�bpP^nl��{+5"M1$�m#y���Pqk�T��N�����J�����hf	ܳ�4���;P��ZN`�Ow^p����V�s��81RÙ���Z"�(y#/��d�h� 1�>�`���]�b�CZw��?����*�ʄ�-9�VtD`�����Xh�In��^T������egRzeY��?d�諝p��>f�3�M����v"��bSl^��ZV��Z���R�	ۆ�4�=�л�2��ȃ���e���P\��ƿ��Wf��Ig��t^[�T�BU}���ዺ�cAM�,C�,����JY��EQk)�o��`ϰ�S�'�S�)|Zw�U��ԕ���7�}�5�����i�<ž�+h��%���)dX��4-<�Z��	�ؿ,���M�vp$#��a���N�~pa��6�kIE8ب���M�l
Ѥ�4�
��@ע�-�f`XII�:F���)kj����K�ƃ�� �f[��N�^H$���ͬ3_T�y���J�T��P�t�np�O~�����_����f$	T�&᥋9�w#�ī~�7?2����H!r�J�eAo�YcfU������O�߯&QQY�al"n�����:�u�	鳵�����:��q jh�t��#�>BM$���կ��;m��,L=����0'=�!�I���� M��)� Z��X&/�c��%�1A$��z�L�JxR9��y���pV�zg� )^~x�i��D<�}N������VF���~����zS�A�����u�L#+J��j,�|��]"���@��#]��3�3�1y	�������є@|�����b}����$,����"�I�_�	�����h�uc����ѣ�m�wf�x����:mNn��,+
��p��$d�&���5�z��L%�jH���K�2!l����uQ��G�|���ר�+���d��^����H�F�ԕ_�ex����[�\jD��O�������(�MlP3^��"y2�3ݘ�*��c�:�[�Xs���;��d��Ǡm\U�=��������0����2�k��/y�]H�j����Ĝ�׵t�5g$�ٌ���b�S����rgS� ��^$�2�aO�]���`����gF�8�:*T�l��Eɀ�a�N����rR��u�ưE!�"�ES���C�F��	�cs�6��1�	�=F�¸�%�������G��X��c��iֿmB!X��яi��yr'��~D]��4�J����cy���C�k̍)�]!5;ar�^�)�_�Tm���* ��q�x�GF {�jC9l7$� ��+��~`�;�`����N� X���q�C�W�GeŊ'�G�@�1*ͥ?S��?�W�[���O@OF&K�&Ԡ�E+X$����/	��/ߞ�q{�4h����#%!�-G'�`�aFzޱ��V��2���o[V��l��yAQ׭��u&�f`��9:l:���)�}
�Ş��rM��dy���A0oj=�sbe�u5@ةbeTg(U0�k�Q&�{̤F�vq2�_b��$��<֖�Y�)>��r�d��تKB}SC���xY��f�9 �'�D˂�0�nV�Y���;t���ml/�4�"�r��U?_�$�㈆`�"zsD��xk��6�%�n�&P��%��Ҙ9��e���+tK"���Hf#�`�6C���(-a�"F6k�0�Af9;�`��BԳA�m�@�:�6�`�e���/l>�9�ʱ��e6FDq�Y>����t�Q.��~YX������}S#6�I�y���E�<D��<�������^e�{�L@2sH᧔n���8�-��I�q���(X.�Oq��h�r�wm~�c����A�8��p�{��V��9WZ�J�B�J�<��arS\=����X���%H����j���	a��<�R��6DpW������DAm!��jbgT����A�hI�U��u�����Xp6�L�q0FW!@���e�JZ�%R
�Y�"�|�*��rJJ�W^=t"�|7���/�Ai$��u0̭2���%8۹=�y��e�G ��r� $u�ZB!�w��1��)	�F��1�Z�jY�`��YC���Z�jƅc�/�:--d�w��[�����U�Y���sz�?��\�����
�#�D"ܤW�:VY�>t�,M���ͯ�8�i+3�ֿ	�ƁYP	[���}D� 2M�w��r���!� q�e�ѡ�2}��*�8ۆ�*��]�#5�B�B-v	K�k5ԓ<���2B�v�ku�l��������ef1����r�ʲ3��U�`SX*�#�t��T�� }5�E����p;{z�j!ҳ��k�D�\�:7lO�UZ������3��0���߽����Y5]-c�5��a<�:1�I�ֶ��t���K|aQS���Ua�\����x�m�7N\��ۀc�����S���0�؀��Vp�p��֞ f��yOJ�=��'�Le���P�`���.�¸l��g�`tR��F�묎��s�k
f��A�e�:�,��07;��>��lQ9�f8ar����h;�����1��1��Yg%p�^���X,��J�s�|��oȺ391En�uX�:	�̡a���j�9V�hɞ�x��̰�;�Z�"�R�T�N|�E(Q*��f��ԛ\�i3,9XL��c�P%45\�� �L�ʄ^"	@oI���i����h+������j@��I:Z���~�1�8Z���|���W��y�p�a"E~��\�� b����0pxl���f��-h�2��$�)�{@0��w����|xD��{l�N�2���z��{R�J�i��ˆ���|�����"�'�<p+�����*���AP8�F� ��$��EU�!�a�z�.�a�l��s$�3	��,�=��`�+kA>Xȱ�S�sw*T�@�²5��
6�O��sjn���A�8�V�GK��̙*5IU](��iĤ]��ꅃf���.�D�T���ذ���^�|�Uj���p��`�#S"��H���9\�R�P.f�7k�Z� y��4�0SB�)�0Qh�� k���A�W�PN5�ǋ�!�.!,��4��w�6
_�^:��6�?i�κ�.�3�Bk� ]�4w4(+�V����+���q��!��ʮr��gNU<x�,�9�J��k���!�/��/������l��X��DM�9��3������m�B��5��~��K	����嫖�*R+4`M��j�/c�Y*�7�^����>Y�s���k���L�'��[���gCk�d
���o��!�^�*�|���oD"��p�f<L���:����!*�i>h%O0/S��xMkɕ�]�=P	[}�袇#���Gx�ɅB��s��&<�ÙA�-#7�C�<��i��ޑI����Ӡ��ud!	?��+�����$��׽d�����w��?\���2k����ǡ��ze��Eϳ_h:o*Yh9�՛�����"#�rK�4�4��W�#�D!�uM�N%f�٥�������A.�x^��+E�[�ڸ�T�6��\݃�?��ݲ0�RCRi�P �#��DJk7��3LG,G]�#f6QJYѦ+������O��5��e�:�:��GS'�wG5��9�~d�7zr����
+��� P���A{�w��U�y=���o=����'�wn�Hb�����9������<0IRg'�z戼�j�2���!U=
1��b�T��[oz7�4�����e�U5^��*�`�^u�<�e��t�"�}�юhf��[��v���BܡX#����,�K7��\�faP�z�S���L{��i?��H�Å��T�T�?��|��R�λd���5�����x�5��͟/���q�e�O�����DmE���N��\`lމy�����)w�ަm
��2�U,\��okK;:�v��w��f���'�Cu��u����o��Z��Ϻ�s=�?�e�ʝ�UQچ�F�h ����2��+�ߣ�P�a���e��F_E�*���T�0�n�1T}&5��H>_�`H}��ʊ��C�>�G��&ޖ���e��XpgH���"-���k�W�.��*JV��g<�<+G��;VH����c�h5�Sf�'\)�&�K��V!U=���V��@e��c����,}'���T��\D1F%qռ���cYg��-V�)�����h|��Z��D�����ꓧ�|q��Ԋ���2A?{�8���vBo�W��N"���?���]~�^�زQ��ݰkJ|%�W�l���0{��4'x\`=�h87��'0�Ra�y���R�73��L�|",������UЧ��9�e����N�{��]�1@��TR�iw�̉�-k��R����d\P��9We~�3��*b�ޓ�x�im�/J������ˣ3����j�L��1�ը%�{��8�t$�^��y��������'�1~>�o�ǲӛ�9���$��ܶ6��� ��=	8i�Y��q�w��"�����8��ÊG����
�2ܶ�v7y�=�"F���&\b�%�(X�X���B�GS��وBoV�vlM� ��	�"*�W	�܎�V����W���%8Ar�����V���I|�}�=�o�,�����.D��1�L��1����5}�#$GEq��*�(�l�NݐZ�UП�����v��UB&1�F��3�U6���};M�D_�E�/�r�@���8���1`6�͐�����ʓCb�G��4����Φm+��3��+�8{?�bXY+��e2�>��0��@��j6� ؼT,B�V�`��$�bW�Bi��t�r�<�bpN��ҁk��BZt�׸����/m��1!�zc�����w��/�D�c��]��xd>��L�V Li�/DW�\��ob���(����1�xJ����
��K�[��Z�-�����*( �������������D��I\��vcθ��7/�q�]#G����+���JP7�K�t���D��a`T�:�	tOYi��DA��o��YM�)+�iW2�uv�r�F6��Z}���gQ]m �>�������k��'�Z�~-r�N�<���J�wrr�u�]���/j�ף�:.���ٞT8JPUb]�`T���J0�i�����B-w`&�1aX4�l
lޕ��?�D&��!,�x2�H���I0���!��njs��/O�^�eG�����s�����π~~-Q��3[�L��4����/5ܖ�/,��5 �����Q�龜���42U����E�S�s��$�z��]������3�s��_��7��mi!%5vT�a�[�}��x{�i����
L�_Y��?%�/B�MH�p��ݚ�BW1g���x�(��� '(4�Y ���xP�K∓
�q}����b`�'Ѩy�HpǸ���5nigH}�2�q �oh�2��]���n��)�6����\Q�atDu<��=B׵�b��O~�����PQ�鸑�$��5��zI��Dnx���Ea�I�M���7���g�;��0����uS�.)y�*nML�۾�k��+\�v��-��C�8��;��:��b�aL*MN�7���l�C�����|��� � 2�4�S�1Ǣ�z��g��
�����n3xV�/��ٰn���9�]sƀs&r����U�v��+�D���_6���Oq����ɢ3ډ�{����K����j2��3�we8�'�����Ç� ��f�X6��?2����#�;燽v��s%�K9V�������,��������j5��i/ݒ�{7Pz�5bו�K��cD�	(�UL�]��xt���k��z���v���U� �����,m��X���N	|Dp�"����i���qC����`��˻��N���%�.�[�s�@h�PJ!�[]��ߘ/��o�იHm�����7XAX�UAϤ�����+I���ѯ7��Pg�ޗõ5���� t�0"�L�^�(	�ғ::
i����bI9�l��qEq�I6��i�]�Mck��Ky���Eg_LE�!G������ ����E�l+��n��y:P*ѭKØ�2N_�fof�r�vȪK��r4Tz�1	C����솛&���۞F�y���O��ɹ�<b�8K�/���8�4P߮�ɧH����N��+p��!�sv�dQߔ�V��|)�p��d�`�¢b6�S���	p!	��q䙱T��ȣ7�m�v�!��p$ڐ��*D8��h��l1��ú��3�6��� ��a?�	-�R���vvˁ�(��,���}�$y3����ߚ�yŲՎf,&�ʉ�	bZ�_E�[(��	��r<��U�7(��(���4��U�晗�;P^���! 2Mٍ��|��!TZP�ޮ��b���j3���mcS�k˪G��R���@�;Y�� �'4�um?@���߳�X��qN�ȡ��TH��*#%�����s��Eݨso���J؛1�P4�w��4-��Cٺ^ޥ
��X�g��Q��vV@��WU}���3�7���4��z��K��=_��Ar��ۘ�����	�����v��v-�>�&���X�,?��
R̬2x�J[�/��5� ��o�F25�'W�ck�&q�9��.��'�ϱ�iU�W)�/��85Tl�c�ÍR��Go��#�>�S��7���e�H���.�J`��ů���vW���ܳM�K]����,�t�(Kq��|w,�%⌲n�gic�i7��vq�{k#{$��w�����b\���i�Ų^���o�u�	^���DaZ��l}�b����LG~���t��1�#E���!"�j{�n��f�F�}���.V�"|x�қS{�%����w�}[�}R�ֻ�ӓ�%d�`��{4^��'̜E**i��r[� �&��t?��H�r�����ՇH�so��ס�m�Ӂ dW~�,���"���ﲵ}�j�r��G�Z�MЭF�e� E�}Ή���Ӯh���H��mr&�A��9�?p=и&[U����Ug2��ig)f��B˹��t^�P9I�*(���4/��}˗�v�~�)FOOޤx�)¢�sb��ʽ��Ƚ��Xs
��(
��P�2α����X\tS�YR ���u��Ÿ�آȌ�T��&ߣ2�ؒ��F �����닀tW������?ކ��h�.�i#
~i/�M��ǜں:荪�*�"���2c��A��w40=�E�)�rD���(i+�.nz�dݭj�4s[7��G�#wr	ɔ2T�Lՙ��Cg�.�[D�D�pv\�¬�0�+�r�0!�b�����|+Y�Ξ;<~���i�q<������ZY�t ��Ĵ�`��0J��<@�r��S-���
a}eU)�C�"1�*��ǵ~O�����̕�@��y� U��n%���y#'x�i�����RU_r�����{����*|(�4�҄��,��zr��F�|��秺C8/�z��o⋭��a魉��e���1&�{�M�Y@���&;Aɸ?!ߏ.�p�_��@A���h��&����T�|J���������q&<���?z�K*/q��N�'��-F���8K�r�H0"\̰}�v]+yQ׼ֱ��U`>�|�U}�ޑ�$�mwR�ㄭQn�(m9!�� �Ù?��F�Z��RwU^�K��<�
��ׂ�:%7�t(ݛE�8�o��%�`bC�9+U���B��}����Q+j��G�Uz�,�a���s|��F�d��T��*� ��iW�x�!O-��m����o;��Y������⸬�&\R��0�)\.D��Oebd���ǩ�v4��@m�??Ĭ{��%Y�)�Z���c�����
��0`zݨzl�N۬vCpOL�}�d쀕�<	��ƻ��"zB�u�s�Ǩ��~��?�n˓`�ں�>��|k3����-$��N��9�Ԡ��N�i�%/��kQ�5��l�"��j��n0�/!�SB���o���6����l�������]]*"x���|c�E�����<��ic�� �g�O��q�_�CKn�� �GL4������J�oy�D��r!���$} ���M:>�!L(�^�b>�ǉ�|�pI��f�G��]	ܫv�5�d?33��e�Bl�ae-8VK�i�>T��](�%ds.cO��)tB�s�1~+�ʮ\ϔ���2U��/�`�9�	
`�^JɅ�K̤i���?SRة\�K�"�NWyٷ�ъm��4��`�G��0I��aѢX~���Q5�fF����oa|��$�Mw�7f����s&���25�(Mr5��$\����7���L�Cm�E�U�d9��^��qܥ\��u�h�fZ`4�U��2��� �ǔ���w1˳b� �ѡmI��;�P4y|1�%I��ų��D�Vf����g�օ�-¢>hr{}H+Eb_�EO�w���=N�p�������^��L�?���q!��!�5���<�愹	}��)�������LД?$&8x�从��K���x�T���e7kA��X`)Ɇ-���|��O@�|B�)G�B�A�0�$'�ӽ��N�5mX�Փc��5����<��R�`wE�u�%gC����Sձ�C�,�������Z���¡u�H�;�U⥴֐�)"����6���!���S�z$�wZ�y�nH�%UyP�D�^45�<̭���PĨ�����b`��@�>�����tTv=N�����~��@
}��SZ:�$^"ԯ!�U���c2��+�j.��2|if��s%����M�?-���?�-�Ӗ:�<L42X]yu��֜i��,�5T�}�2�VO˼!��E�Jᴛ�
�ê�,iQ8[��D�K��c�k��8�62*�O8t_�#��p7�&�f5o$�2S�~�x"�K����̠�py�Ő^�s�;�._]��~k�^> 2sh|YE���t�//��%�$���ο̎����D��15����u���'��Ѡ�N�^��j��"5�j�4�t��ڀ��[�hM*O�d�ڑ�I+�m�0���9�܃��n���S2i�9ձ0MBɐ"���5���߈�D^wH�[֖�q���"��y�q���NM���xX�@�QS��`f��f,����T$���t����Z�c@�n��R�z|C��r���+�N�H��T�`ꅅ��k�nI��	��]ֈST��o�jD��ԍF���m�s�zk<�UΘ��}�&���^�qS+CLl4���]ך[��$��#� K�p�XTя���&��� �k�����O����"j�N򹤚�~�|�
��,�����#y��K�hu}�������:���U��=�z]ǮtF�i�N��N�7��������Q��i�z�~2�J�(Ĝ��?S:���b��K����~{[bb�*���<?P��u�P:ݔ�!�I���5����L���!��:b�-�<ʙ�Jj���և�l���q$�i�,�����wibΧP�� ��Lw��Rz�2�s�'Hrv��jio�_��[���W����#��,N���#��9k�"�����qs�4ZY�-�/�bn��}�Yoe�7�d<i��m�gܼ���&����Y��"RXT�:��fZ	 "������U�!Ĝc��c!���6���1�0(��M>��d�N�u{�Hz���{h�S2w2����Di�S9f8+���C�*����GF�}Z�[J�����z�s�/ws�`H�;��8�[�lCMă��C��x-ErϹ�˂ŦhA{�J�>N�0�M�x���X\���w��*���R�����$���jz+�6M,���-j.f�\0ڿ	�Oe.���<ѿ'CN|C��u�K�=��֬��(^T�&�Z0$;��ܒ��ыf�1%��!���4Y���։Zg궀��pw�T(�(}M2Ao�Z$"Y��2�C�s,�} y��.~��f��rb��	.N;�=��H	ݝ4���Z*�uрB�ԥ�'gx{U�6�cr�F7�]�����&q�SsS�X/Mލd\�D����j�1æ�P�P��
{6��N�P��K�c��ӯ~�L���R�[J�R�k��Aj�
��X-a�����5�*6&�E��ag����D/ۉ䘼*Lq�k�#
������W�o�~>������^�FrMб�5#t�OÒ�Ƿ�Lg���;���[62�����~��68bwu�ItV�l�K�� IE'6Q�|�[P~,�u�O��2�ݘ�I8(T�ryOG��G���8T�O�څeR�eż�����=?α��*m]��57b�ΆT
�ɦ,�KՅ.����ݩ�}����"�B!�^��=i�[�Im��e��u#=~.�k�O�S熔~�\>��E<���`���4ZWe�)������i͵T��.�CI�@��A�㳯^�M�.���s�P�[-d��bL�J��s���3|��E�@18N`p���G�����X�����-��k�@e�ҚY��=c���f�0�>��8�|�	�0��^�-�3:���W��8;�lNi�gR/6>K�ܔ�}d�T�Q�}�r�J~4\�����P�����@�Ay�`f�add\)b���'�e(3�;Yi0�(
�Jvl�yX~���
�6��ߦG�&x�a��Ʋ��9ۿD`� XX�����`�������t�WLvW�futj	�m	�����w	X�9R�6���Ad�W��>%H�\�!a��ˣ��'�}���18��̶`u	��W���J0�X0W��H�,<��LNS�-��(�n�66,�km��j Ȳ�n�����;�3�P:?����w�r�����Q{flN�W�%g�'O�gD<KUx��=�;Շ^Ga��NДH�s,��n���@P�-��|���l�s��[Y^���׽��M��Y}���Y��!޵j,O���B�{'�"�	׻�}�w�П\|y8�G,T�E#91Q�IU|2UС;�݂)X�k�i(�?&�8��ӆo�ՙ]ER=6���F���w�	�Aa�8�%oN����g�V�J��ug\]s�+0L��<�$���g��SnsC�4i��{�mx,���*p�M��ghk��5ʀZ�$���h��ᬈ۹P�k�7��� �g�@փ1O�MڦY}�F=����Ⱥƈ�-=��^�ty�l�H��%ˉ�ϓ*�cA�&;2����G�Y�����m�-GLS���>;]�[;��P��1����(^�C������|���zac>e�m�$���z����3[I��8\_J�C�<�O�]㨫�s�8�t5���O񊢢�y)�ˑk�-_�u�U�ށ���}[V!�֚	�t�I��V���,���aNݺc_�6�n:v�>X��jǿ?��0�V��W�rĈ�O���7oY�X��?m��f������������@{͉|�v�U�iMO�Md$�CC�D86��eĶ\��{/?��Rx]�<��jO�e����C����2� 37>ì�R*��3��F
�f�qI/�k�
�:Y�˾Ѷ��PM���३��{	n�#n������m(���V�d<��~�]~l�'�z���X�YNY��!�G��s����5���(���A�:��s��>1O@�1	�V~�<��y)��kA������zm�R|3�nc��G���k��ױ�4�ii���=k�9����������G?n�
�eʳ���� tV
��Ǧ;��^�F���D�4=����3�?�x�>�����\�~���FH7v���y���KqL8�6g��-gXi껫�>��=͒��E>�dFn��a�4��3����Q7��8ޤtW<n�5C�ѐM@�]�T�s�ih.*X!S�7����#{�s��%���h�)��Pd^"����i1 G���xy���x����7k}ʫ�lY@��v�H�М����!D�XB �q��]��p]���,6�{�e��2��1ک��ht���W�>�ޜ��q�:�Y�Z��\H#zm.�?��Wd����LVC� *�cZ��@<���tr�F���2`��/�|�b��y����6K<߆:���U��?S:��t������=��
��M�Y������%W?�,��c}�Xs�C�3���"����	ӻAͶ�&�[\@��U�$
�<���\��������K_X������LxO[p�<U	�\�JZQ2�����/��g-}L3����h��Np�-7K��j�����3����=��oC�Y�o��ɵ'�}�]ڻ�Gv����c��x\)��zo����/�G�fb^�ܩ�9����"�W��'JycBM�O��s!�(�߃����)~�������7��I������]68����\�4�@%.�����@]����M��r�H3�d�\k{�>�g*�=atv�o��M��u�T��e
L{\_��-ؿZ�jNhΰ{��VZ�f	)}���Fs��JW���@��4ԣ���*f�s㑗|vǺGj��PO��ǡ�Liw�*ԓ��dR�ҝo����� �C��|aG���-;��ڞ��z�G�4�3�N�n��7�z8#��z�?����4�	��@x��JԴ����pFg��#JA~m���� ~�?qz�Sڝ��c�k=6�}M�T3��ń+�������P��!����t�o��N��z@6J���u�_���0�g�C�B]���[9|Pw����3۝�z~ö�9����D4�]e�t��)?���W�T]��ĝ���n��^V��Rm&[����˹���r֔��j��R���~͸UK�)�$+����Le�⏡+<.��rN��FLqG�<��KI���Xꥉ�ǻI,ѯ�b��#*�"D!�fٟ��N4�<{�'��$�֍N��� K�"�T���8/�U���>D;IS���-&�����m�3+��F	�	 �x���`�.50��+�ِ�5hj3�oU���
�X��,CBۙ8*�/�&��Y}�ABzE�2�#wx7`J�@Ō2�+��)�cw7�����l��^�QR:u�"�|�vdX�o�,�F��k�Y�2H�i�.�������6�,���`����z�
C9,��/�7_�*f˿k^�
?��J7�b�I]���.@Nf�'�����Y�{n<R�P��0ZR�Vo󌐒	���oc�>՟J�҂j�H�����#�UWǓ!���Z��=���-R��c�Ϳ����Ɩz�[�Yd$f�R���p��A�.Rk{p<��A�f�tH�f�hd�y�b�3���َ���ڢ*�[fY��sw^0�5^3��>2��|ɕ���6��<L� =�߱wa��w�eCnd��X���%��R%�)��1nfU���r�t�$2�O�h��q����U��_?�W���i�g8�0�Ր �z�F����&��;�Z�!���M����4�8�NR�Q�:�!/�	۵�1u��*3��5K��r	�&��cln��F�~F騚[5�,��X�M��6�1�]<��8�/N4��P7o	c����<C,G��t����?�����r�b���ѐ���VCm�R�K�7"�G�+�2�Z��ǟ����`�㌨@t�p^8�ې�1�%�HG<�^�/giW�G����K���j��ˡ]��oVp��q�Ν�̮܋��l�H�T����W��Ɨy���H�s{��>�t�R��k��r��ɖ�"=�� ��ݰ��Qi�2c���d_ʨ5y�.�XBW#��P�0ĮU> P]x��`��	!�\�$z�y;l@�[:C�6�bzw��9P����t�d�CR�M�^H^l�ͷ���bGh����6���E��ܢp~x�;���A��­	sr+�vgv�"���cf����#���Ⱥi�O�>�Z���U�hk���;�'��1T�S'bN�^ۤ#�����)z*¶O�z�J�ߌ��$�������w�2 "�*����/��������|fs�2�%���m�.���G������2BO��aҁ��AJ���c�Y_��	f�M������\.� �#�Ȩ��ϱx5t�bS�GG�����v��^�[���8�N[�w��F�B֞��n����o�{���Hr��w�s���7j	L�Ɍ#��Vr$���~�+���5����=�q��w� I6�`i����f�n�<�^	�Y���_DK�������?xc���%�r-����-�n����~��!��ϖ:���|$w=�Uq��'��@*WLZ�hN������>ܰ/6⮆g�1��q����~����sp�i��za,����\O��i������Q7+IH��:�] �%*�*n����� Yph�WD4@�˴;�o�vP��Zj�˻� ����ˇ��V��,t�t�Ez�6��.�����j���������.�D+�L�I#�%1�&�]�����l#�z�U�; +�/>払<,�]���~�29���05 �N��I�I����8g���n꛺T�����O�v�PѦ����U�ن�V�dc,�#�I�B����o��
��͠���rCU�>g!�p�0�P���6�J�R6i��(�J�:�K���s�s�P��� o���@/x��Sɝ�}ck��v�g��n��_bgg�6HT�3�!��BPإ"�/��\o�â��	��]��O�>���xN�D��gu|���vL��F�7����'|}_�g+�I��	֧L�>D醒��8t�pT�6Ǚ���g"� �N9 �;:9b���t�{ �煽j�
[za��4�^BU���qߥ���K�J�F\�[�zwM�zHX6*َ�q�م��E(����H75�j57c��&�S��C۪yFN
�O���l�O��"p"�l�'��wD���ګ�\h���m6~��,Ŷ-<����J�gx�[����x�E�v*�S2(,����kw}&[Ȥ&�FV�7��������b|R����1?�i�{�u��&8T�����t���[}G���T�5vl��?�9v��[�±"�0�bZNB�yd�M,�􊭻��ܔ�R�&!��ܜ��/g�ߖ��WHژ�˂��[]��Ԙ{����O畹�ɒwF�_a�k�sy��t_����̙�;�ǃ��o^�gd��堂��+z��3����SU��z�~���>�A#�=:��MG��W+���Nhإ#�S���,{�W����p^�$#/]C���hF�E���;U��B��4GI~\�lQy��I�>���T�zܗ�#ȯ��H��j����Pyn�FWe�f�k��q=��.����*
�"��sKH�GC4�$�ز�v����~u�C�$-����֩E��l���FFG��
T�za��°&�~�yʜ��iR�1ǀ��)�sh`����k'\p.�)��x&�ĉ�L(V��.��,���?ĥ����R�^��]s$��qҏ[�4��,adR���?�`ͤW����j���Al8-z;а�o���\_���lQeb�]�q�4ïU����-� m_�|s�"S a�2n�6{��+��@��_��W_(�1��2x Z���S]NY󿼠45���ܥ����'���e����a���٥n)�uB��_�@�ƚe�A�#�x���H�i��؍��!�-���:҈׳"���qY?6��Yn@=����K���2�|��'To�&#U@?wB`>~�91��>�~AVD���R�b�j��!��l��p��~�\��kA����)�[x{����sy��S���`yYC�����9�4Q��k#�ܥ'E��G�n���i�Ed��̔.�����|w�0wLLb�X���]�2�ZMw��_�,Qȶ�νb͂cPTێp�D�i:�Rsp�h�T8�#�f�hV�$�l��Y�>��CNN;Q��&G�6�]���#QQg��邀R�����-6n�+�����r����[!N=�A��DwcX�`�������kEJ�\�[ہOM�� ��-�2h�c����R��|lEj�*
�!>p�7���ڑ���|�w�W��K)�v�����W׆�)���]��Qz�Z'�|��Z�i���i�1��!.���%/⟒`!p�� ��/,��n�n��*�7����v'��/ ��j����.\]?�}B��y��N���T�j!o��Fҁc�Bh���ߵ�+�Wtb-s@�؇���9��٢�ۙ��V	]CF��(�)2מ��Ο�'��4߃/-`*�+J�)��~�����>�����8mhWrMIW�eN*g�|T�J�ZCT����U�"W�>d�é�Oؼ�|S��$,��+3�aF���O�' ��Ê������h\7��쇕�hj�)���s��ӿ��o�MM?A.���w�������b�Ɲ9��;�f;6#��j/��
����;M٫p�S��Şp\g?�Je�q!�A�k>(����\��O����1-X�1O=M`�_>`�[���F�E��L��Z=K���k��s{t�n�����9�}�����
�D?�f�ώO�BU<	 �h�F)���j�P��T$j��-�UF=%Z��"��X��;��^ɻ��6<�X�n�M�Ġʙ�TI��'E��$���X��F����OT�5�ry�� ŀdX`�hG��:1��3+���w �}�$��6u�g�^ꌅ����7����|ձq�Z�Os��!��*{&�>*y�LQ��lN)�ԧ`���>@ӗ9�~v��1i4"�E"/i�3wHc�!��\��kDu��$�8i����\�_~� 5��~��3w�C�ջ��~�����]���b�4�/6+��#��YְYH�qh�T�D�1��N<ӝ��d`i�4���ز��A��u��0��K���<��k�ȇ�9� "�X�q�A>��3*<�w��L���7ђ2�����K�k
����ڊ�[��hCo��Q���A�z���.}Lujn
6��0��m+��;y�ɡ���b8�#��܊`ɤ_ ̹F+_�BU�Ԯ��~ro"����*�@w�q��Pj�k�1o�A����eW6���4���(�(r<��?�A:����	��m��=������l;�=�})X :���ś�o�4��@��˚�1������Y�����X�?�@��Y�:��`bM@~>Y��,&�L})o+؃��E�C�z���H���(̬���ҹzS�{�u=bX�AJjX�-��H�t5j!C��3�3+�n�b�_-/̳�=�پ�;+:�
%����{��}
�?�c^]�b]V�F�>�Q�9C�u���X��6�<�y�7�����N,�~3f��}^g�&_��J�Z��x��Fk��1e�A	z�ޜ8�S=��A�=,��>��_�`~��5�� ����:�,�e�^���k@���
S>=I���5� fFh����3^Ε��
N��X��a�-�[�-L��6�Mf���Y9 �J������?)�l�֎PE�g�+*����{�}���&6�Ɵ>;���c�S�����?SȶH_*R���-2���r� ӯk��^]._"pt��>r��w0�e�W�^��-A7_���|��;���tT�>��o.��;��=��Z�mi%L�:���q^����S�V�$�|p�^jǂX��q��Vl@.G�L�f���u?(מc���e�
�m݁?jne���ݯ��b=��2D-|	�Ɣn��a��]��%݆�v�,���{hD�|���������G�"<"��zA��*{�w�.&�ٖ]օ+�Mo�׾�u�[���,9�C>!ǰK�&Y ��x컲���2�|PSX�L҄>&���
-b�^p���W���Ώ ������1�����5��h/v6{��ĐPS��������������cS��Ls��3�t����*E�C�S:�����YU��
���5�Ծ��b(���C�&�����\��>\>�c��Њ	0�MZ��(�A��:�Ա�.@jy��_���,��_��3J�O�Ql�_�&U�dND-���J�tLJB��I-�-�|�&/����G��8��	'�*�L[ޣ��܏��:oX�$����F����Y��"\G�T�n%��i�bv����H�g��ȥ��j��~]DQǞd�T���&���O4I�MՁH�6̎ �Y�p��uv�k�y��+��jsV�c��m�`y��)p��o�ʩ͍����,��s|���gކu���-�ƹHn�"�G`_>f_^/��u�免�����_VO����.%r^\Cf�db˻��Œ_"��,<�>8�����o���6�~K6ĉ�/�R��/�VW���#�
�a�h#��xi�����������܊ѽ������[�7��A��CЏ�o�=���I��u�|2x`~�K�剃hf�a1��%w��y�]=�����Y��*�w�/��Q^�}�J�CБ�9�J�s#º�62���ѭ/��^�"C�(:"��\�~�^L���w�Nz߈jQ��	ؕx�#¶�|���� �j\��pj m~@��.ܗW�cX�37@�����$�U� jcD��{�5��D򖭥�Z6��#�q7������0D���[HX��	���VX��A�#0��C���Ѿ��6R�SI�%����ޛ�MKqW�z�郴� �i��Q=������@$���?@�ka6��0�EO���������.C�HG�{�Qǀ"^�O���CL�5��v�Kf.p���F
dn���hV��۹����7�|����j)q2|��������_��h�Ǟm��'D�;9����9߃O(JF�5�(e��hx ��b�FG�<�c���	ksi�G�v��dN��#���F�#�;�`m�ZPB�h� `�m�n�H�̸��3�'�2��9xb=�������;f��;��eu���O��r ��ACa�b14dY��S�a�6`L9��SÓ0.h�yˠ�H��Q�!�U�a�sXV)ݷ,���ѣ�6s)׍�z�G;]�9��M�_�8���|R�cT�r�ԧ��\�Pz����\���2՟^�ތ�E�����]��������]��˗0l��V�q3}�{p(�ϛ�O���e��39`�J���Iy��W�+}&�,"�,�U�Q���* x lV�܁�G���YYI�G#�w߸�.�����6UYy_:�cU�x�{A�h;�=�5���-c�+v[Ɋ��Ǥ����m�~c�qP��ʐ�X��sn"�/����s����)NgW�1�Б�]>ͧbF�X�{���Qx�?���إ.�9L�	`�׮�n���s8���S�Y<֦�L,ˊ�Dʔ�}�0Q�%>BĵńL�s��;�3o�����$���D�	�:�F:ϼ����<Gt/v}D,`;z�#o[��'10�li/�y]^��%�����Ә��ݹ�;ݮ����X�'��^�l|,�e������)���k�O�q\<��G�$_�d�R7��fgt�&a��8u��H�
���N������)L	e��d7��� d��Z�8W����R3Y���W��{��#����������|B{��!��	1���5?{n&�N�*l�=�X9cBriPj��u���g�T�Q�U��,(%���^#��nY���^?��o��j����56ԝ����L��^tDpփS`���9�6�{�@��L⳷w�����* =B-�ӯ��U�/����U �|O��z�����V��hV��������@�b�|��x�ƈs
{�1�R6;�U���3�Ֆ�j��O7�g�p�W5��N�1O�v��V̌�H��_<�ӋD�Z�� 8�x�
�Ƹ���\��a����|�=
���0O;�,!�9���s����CS��>���4[�!�ՑfH˿� ���V(�/1H���>(k�����XIl|7�ڧ'�F��~\���$�&��b7,��=!lb�=�dw�̠ucU�î/��n"�9a�'��U_N~m�8�޽e���-8�
�aR)��A�6���?g��j�J �+��fD���L�����0v���]��J�w�ۼS��l�[��تq�G�X$�+*����	��=�����[s�`Zͥ�|Bٶ8hs��_٨#X�e��&8����Y���8�`(��
��Z�R�>��)��nF�jwj��s>^aؕ��2��A�H�^|�:��c7(\Dp�؂���E��Sۍ<��5�A���a/�$�L�A�夶����>,�q;Z�/��2I���*�P�a#i�V%�&�2c4��!Ի/x��y�)�p�ǐ}��K�J���'4�t,C0B�s6˝_�~9lD����@��ls����e�Q�AH�S/kV�~��H�Z������S֭�&�l���VҴ����,yy$�����80� ��.����	�݇	pyn�-������Z�f�vRf3�\�Xe��a���0�%��S|Aս1ȭ����=R�<� �u������fM�A��p2	�stk�YQ�z�u?3�ѫ�4<!l����a�V���I�ۥ�ic��v���|H���\2k+�6~]&}��UKj��� �Tu*�1��a8�CƧ]��H���+V/�|@�9p�h载L���~H_��[gu��[�p+)��[2!jJ�[�p�kU�IN�v/��nO�~�$(X3_���C�@PO������êg/���Aܦ��?J�x��ۣA1�������������]QJcs}�M���� ��[�,Q���9LK
�L
.ה9���m=,V	C���Y�/j+�8�+v����\O � ��ӡI���PJ@fl���S�E҅ �H�t�������p�������ݼ�ҟ0�ْt�I�=S�
*�=0�2|�p`;r�޼U�	י��8���g�CWy5�\�2"���s���^��5�2ݱ���0��g����4b}艰�֦9P;4�h6Q���u%�1S6�Ҙ<>}qR5,�Ry�t����r���!�Z��MQs�L��A����j� ��CÇ"U�	��e��]�=>O�63_��~��?i9��S_k������1��$����\@�a3D�WL�P��̎b6��P�h���,���n�j�O|s?xq����
���SC�h����qp���c�K�W�/�3-��������!'�D8"��[YW����ഹ#M`����+wt�KQ��h����L1^�FCD/eI
�4�����o+�U���D�f��uf'r�l���)	��sm�n�gM�}W�q�j���cDc��6&@�Wچ���!u�ʏ�}�}#�����-��aEi������q���M幭"�ټ��� b��M�7gCK�&��!g�>!,ؕ�AU��a�׎O�g5ÔYT�Fܫ�6t��#�&��'F3{��IP ��,>(��.z�ڊ�_��EcF�ݬi�w�OhQ}�ڪW�,���t���	��u��_%֩2�����ABD�~��c�i6�	�G���'ia�p/"p9b���7���
`����Qc�5r�b��~�~����'?|��[��J'��SmL?��08��gy��]i�>�����ag�B\�\��HW��A�n%ϋ�	�v�����>�!�IQ`q��m�J���}!2^g�8�]L���Oټ���_����˪=ii�SK'� �^���C�=�a�H���ѐ�G�F��(��w�y�؈�/a3_�����+P���$t�[0
�����F���(�(���Ҏ����s?�d��E��c�8�6Џ��
�̖��e���_�u���)T��ߩCJ�LB��dǽ�!��a�c����P	R�5��]̴�'�j�QP�}FŕI��D�m��ӑ��|d������)���e=LpN(��Zu� ���Iz��a��酾-o���Ԉt��c���8�|�Oċ�hnoaW�0Sx�z�ɗ�`5��i�5THʣ!��j�__?���F��g�����w���QR\	x� �H��N�I��U�x��< o2���uW� �థ���?�=�n�@��ۧ{X�����?�]�_sLΖX�M>�?��ۦ�K��`��Y�E�P��n� ֭�R��=x;E�ͪ���fR��	T�U�n*{�nj�E�D��"RTw�<�뵍r�m!�U����R3Q<��>AM��v15�kI�R��B��F���me�av$4:��.E9��K
9g>�C���=�oO���j��7O/��o}iƟr��VRm�{�Y_ĠN^$-f�f��V�Η
�Q�n`�Af-���$�>�a��b��������Y$?�w6$ZU6b�(B�	��b?�`3�-X�9��T����69�v?[��^��H5�{~܉B ��F�eS�!�p�����(E�!��7'M4�s���+!5,o!ʯ�?��X�I�(͝��ɟ=��I�K��	3�&]��X�[������֬���ϭY<�<�q��f���>�4kc���;+pR�4��Rls^�Չ�I���=�)�ȹN�3��5�+��9G���Ԧ�%�SĪZlQw;=�0*��O�ig�Avx^NG���M4�t���9p�8�e�����+���� -�"��>=�L�<u;K2��<(��������
������n�T�'��|b~���Tm�Ȼ!��Vt��dF1~�}0�I�Lv�v�)	[��=�F�f/���J� �B~Ǉ�����0Ї������N�u�/�øݻt2h�_�i�#����cU�"�����A`V�܅F����3ײr�@���{�frT�&w:��!z��/�``7�Qe����v�� �CE��u�EȣSz;r6�^?��d���Gf�z�@�{�erN���'��柄��=��qtm�<��phr������)ˬ-���O�;�'/#r�F#ҽ��6��eg����b{T-�'ˀv� I@���И�;�e�M�$�B��]h-���j��}��R!���#D����T�����֟X�|�^=v����1zR{@��9Э�jÐ}s:�V��$[�~"� i�|r��@���mK�-C9j�8¶R��>�_2�U�F-U��y�v�:H^��_Z��{a�
\��t�H���ZR�~IM�7��_Kgh�-2+������XW~�7û�1�7X�Z��J0��&|�̠���s����u��1��h(lѪ5@��&E���A'�`eT�N��p�(pS�����I,Z��<��Bj�a�w��Z$T��j�W���3�-�@&��^u�s}p�Zc�Y��2�(��ʄţ��>tJЇ�H�%U ]p���Hv��D0Oy�-T��{&ek���=^nAߩ��# �(wQ;
m����a�ѻ�A�	&V ����5T�&#솲�͎��1焹��0=���4�2���`%l�Q����������tS�I��+��wq��4Θ��w�t����=%�W�49��T�Q �yg֦Y)����/����o�_����a��\�m0��9&Y����IPk�Ftg'}���=�C�g��v�����Y��]��:q�L��}iSW��:��*�%VSxiܬ�AMp�Ә(9	?`IL��``�=
�L��
�n��"D�f7�щ�����Z!���9Pԟ�]���=�.��s���]�gL��!�������(T*�榗˗�E�!��TA���9/s�_M3W��d��U�Iu��_�H�.#��gIثg �kC@����u롙4�@w�����;v��!^�fi4 �2����a�1��Q�+y/��o4��`�i��Sˇl�ٸ�&q��p�Cv ��gp�~��9��vW�ԩ]�L?�I.��1��<�;Pܯ+�|,M���-!�@C���%ب���ΝuJ�h��F��Ƨm��zf���+
�l\tp�+:�\վ]t0�X�Ao\�I8��Q�\�6S�c���L�{���֒q��&7V�Ɠ���`6��+1%W]d�{�O&7m�G5���1���wY�彘Q����+��QZ~Re
�*̦
�^�t,1���M�)��z��*�q���~� V	�JK��pQ�Wi ʛs� >3�� ;C���
w|����Y-�u�R�wU������d���8zD��ѹo�9��>�|�����*I��ovX��n�g�M�MVQi*@�4=f��"�/\���i�g�π��������Ta vW+�!���W�f!�&����4�\��n�E�nN���pj��M�������Q��]]Nrf�|�Y��3�h�LJ6iBha���DW���1�w����vy��\�;�<���r�c�h~G(�� �qށұP �,n5�J��%W������@QdHF�U��v<����)��?�ӑ1dk	Y�lN�ſœ�XlR��������1^U�̓_���G\'��Y]�����Q�&)*��pO	���}���F���z�պ���8��t��S=�"��ŹA�Z}̈EK!¡-?me@DV}/����&��踠7�����:�rh����A����f`z���Yo����]�$_�ԛ���hRwFk�y��v�!$Ʌ����aw�HJ�M���D��Ō���T��W���I�K�*� 񠢌�b�H����ޜ�<�Yj/~��x�S,X��	S�ڽU���!�]4Ņ&��rsG��J�m����������ZJ<�-����X���(����obsL�v�L������]�˸U�>����tdU}��� �RddZL�$���w�l�K����],Q�����Ǔ�9w���F���T���Y4u���Y�*aZ!�� �}�v�7IQ�N>��:�"��1�-YV�6¥�&	"�aʧ�w���RY<B�������`_0�Y�fd�߹зRգkآ��m���&,ߩ�CL���Z������&%~l(�`(/��+�C�N	�o�����CF���1`D&�%G�	��_�f{1���R7�E�;��3�
V�z�|,���!=[�I,9��$I�N�����(8��^�٩c1�{�)�b��_�����:���O�[���Q�wzy�'�g�*^���0/4T�OI�����nOஂݓPsf�veE1?��W���,��f���sr��"����[�w�əپa����>�%B��gA"��qqFN�d�{���M+�J�<ɥ4�z��D����4�tT�a�`��J(��%7'nCu]��%��B��e~�H��>��2�s�� ��A̴ bi!��4������,d"T�i
�f�u�9��nw/	;�L�	��TO���WЍO��"֠���s ��K�i�Lнp ��NG�+c0���wRa�y�ܞz�S�l�n9��Lf#�YX�"��n�D�4�H��1^�B�"6���z��2��As�>>�2k��wV ���ś�Ġ^<\3o<�ޭؑ�/���`�&��2�52L[x@~��,��q�A&��³l�!ii��3��1^=٠"���������}6�.��>�3�����n��b��r�^���(�3svM��a�����wa	�NH�P��� )���s�h�`�k7�>�{�)�*�=�ޟ`d@C��� ��r�i�������Fǣ<�S�&m�(�Sv�*z=i�x��L�ģ�u�p7U�i�p�"	3�@j 	�R�/ ق�9�	���_r`�NA�?�9�}�9s��?�
�Q�#0�D����T%J�<�n��!:���E)��A\p��}3�Z�Lx�����&L�0��I�~�{R͆A1�����M�/1�����z������9y�,`��u.�Rh�/�%8�8��M"������Z4�f�h߂~��� (+r�y�`���'��=%�.�X�|s�\Y>[�L�Zg�,t����	lPk���p)J��fG����t�U�k��(�~�!�ډ�%'s�F3�8&Q�����z�m��.���s'%{�餯{S;u�P�m{,\QO©�[��d�� ��r��X�̏9Fe���Ĕ�&�iV��]�������'��1�ݱ�k���ױ8^�З�Ļ:AvwJ�ԯ�ӿ�OO��sO]�j���{z3g�"��0�Vʉ'Sg�5��^��9����S���D˹�w��.�7����e���K�˅�x}u#��J�nr�;��ұ���^i�D���NTKkm5vGnc���kg���g'��,���V����<"X�?/)k����Ly�_=�DFe���,��i�i�����n��H�ګ��/�����v=�� ˼��t�'D��/�_�Q�g�K{e"2�Q�����`T ��+�O��ӭ$f�}�X�msM;�[2��_�x���񬽊���/k�����F1��a�&�:O���s�wc�G��`��6o��'Q���c;e.�ه?C'`Ӡ�,�Rq4!Tˆ���v�N�\�)��1$Y�y��q���f6P���Q������=�&^*���/G�2�e:���LV/)�������/�U�7P=f���(I-�q��VbE�7N>��n$��8�.�-^� �=�h��Y� r(�}y�2��U-����1�c��+��>��h��z�X&3~��s,�l��6���/��ݶ�� ����&J����dx��vC~㑆�9��h�<���l���*S9mq���Uon1��t����Π�C@hW�u/���;x�.�9�x�v���L�����+��c����}�R�����߳��Yo�aWrO�P!�El�(��
����t���Wݞb1����ZoG�$}w�9K{)u����J~��`v�	Cuu�X�ӥ�ҜU[6�L��n�PD7c�y��$�KG����W�mҜ������Α��L� >��i���՗���Ėt��P��qwz��\+hI��*� �a�h�;��>f�֠�H�@Q�J� u	G�����R�6��_.w����G�޿)�h�2OQi:�=��j��A����)�/0J
��
^�75�Lڳ�F٥G�s3C �H�G�7�9f,X"^0�e�铮N"�FNPpܧ��ob@�X����H�9��x��_�
���W�|Iġ'X������U��/�k���0ȊѪ�0w�DD	���!6�,��b�v�U��B�O�	��T�ZDf��k9O��jw+5�Bt)��Ɲ�,D���uǚa��Qן��?Iѭ]q�9pBVR3�A��]��Ȯ�M�n��a��38�ğu3v5�2��@5���е«��|	}T��� ݨ. ڶ�uH�}D韽�e��:�)NزJQ�Y�ؤp���S�qX�&j�fg<�RFNP�3��S�G �(�|�u=�A̙cչ�S�${�b�J)��}����]�	,���*��q�!�q�7�{�ΚY���|?X'��+�B�PLQ%(8`����`�L`�k\0h
Z}
���.�v�$��a�����h����p��7��@GI�(A^#��TmR�h�� �Ƞʖ��+�>��[8�z�Sg&iy�Ǝ��-5���z�A���V��ͻ�BU�����j@8x� !�"Ok��F�1F��!��U�$�N�� ���P� `�~dt���
w��]씾�D�<�(x6~U@I�:m���������OX��P�5m��ӗEH8.���dQ2���k�t�uK�Sb�R�{@��F��Q�1R��4�w4]�}��/g�jQ����	\��W�^���pC���fQj��։k��TТ׋���I���{6��UF�yYB �)�C�����I�g��7�{��f�	;���9�5�]W���,7e��$�ng�q��f�ݷ�eo,�U`e"��uL��i^�ą��q�'m����֨�4,/��	�τ��k�r�`�B
���>sBN�?,/�X����/���Mr���I��r2�T�"��v�RǠ��Fm�}�ЛJ"�I�����?hVhy�F�>P̋�)���Ͽ����Lň��}��y��4�
����b�r�������$MI�Qi��c�~S�t'��%��U�jH9�Ç�5��!\��
�X�����,ۥn����ܲ���U�N�G�'p��d�3>��Fi� 	�k+�^��(��Q�a{y��B;Z]ͥ�ؿՃ��l}�u=f_[~G ����ч/i��A�%���,[)��TCV����a�RHpf0�%�������U��n	��س��U��1j�ۨy��"@�-Er�[�V�k2�$.g��0�g�dȕgFM5fPƇ2��סP\($<-��tm�'�L�ڢ��g·DV�ฑ��+�H�>SZ���U�j��0R���AVM�9�VԝKר(m�^?>_s�2j�/@��o*��[��L�I����3�Д�/6zc�ɞ��D�Q�u^�B�N_�f�A�'�%r>~��sN'?A<�w�L�_�Q��r�\A
7Ь?�y}9���N=���U��d�Ϗ<�م�7�oh3&~�Ҧ��9۱��<y�/�A%��C͢��f��W="©A8�ӷޕa7W�o����L���K�_ʐ[�Ջ�5˗qvk�E�x	��l�P�����g�A�ez�JO�J7��g�N\)ˊU�>XS�ye�Ƣ���|s�~lu_�C�LP��H�+�`��T�h�z���.q �Ѹ�:T�O�N�v}J;9�?[0�$ynü�<P��_������M��RMI���t�'i�΍GK{��o����e��Z�ʏ�XW}S��-���Պ��n�b��T�F\.��y�Ir ��ĈwY�#3�7~^�=����bk�e��B�w)Zk��d��ǖ�zg���P�[����!_�hG1��'D�̚p�@UV�NB�zs�����v�^�<N��&3g�^7�_iGw3�p�T��Om��,��xD{����Ų�5��m�_��o�ܪ[�{(n���J�`S��@2��c�o��X��]%)��?G��//���񪽲%���	� fΓ����
G�{'n����-��Ζ�r:L�T(S�`tUh.����I�wk�#��k��r�ܟ�w0ש�&�e�]Sb�m瞱A�w]�_@kw�x'R"<� }q�Si���*qp�����p��A��aty5c%���F��^��3��P�R s��m����}�A��	�g߷և����&�9�c���eSR��;b=c7=����C��ߴNeȼv_b`H���6/۷J����}������Ky]
�+$��I?;��+�8���Ջ�)����]
�C����9����J�2Q��>�5���4ۊ�n��e�|9�U�m�Qr���G��/�Y���u	չ��jiu��¹^�/�sa�r>�o;��6:����I(���Ѧ�g�WRSf��kX"���,C���7lU�~�G��y��*�?�laV�ݨ�i�GK`GP�� ��ʎ]�z��U=�еA'(*ԓU��<=ٔ� �����nfQ�_��B��i ��ݿ�v�M/ڪ�r�*��56�Do�N���B����]7F5�*^�z/}����%Wx���yN����H�{�Kq�F��i�C�����q�B�|�:�˛�אM"'Uh����BR}h��]
��.�m?	I�<��H��;��F�(�R �Ȝ���\?���ɲf�V��T��?�~�{���	E��g6CT��<�Q���Yd�NCMgO��	φRW:`�� ��dTK0��{��y�;NI]X6S*��[�-���.���� Rb����v|���V�:���ɉ�2��S�{��_"j�9:;9�E�M�<�>��������蘫�rN���k�dwW�AXr!JGD�z��J�����uS��HRѓ� ��J�*���(��0�>s��/H�.Y9+�P�/�k�Y��;c�� �Ṉ<]���{��E�c�ș������A����D_�XKӘ6.Kvj��~� �A�Y�|2������0.�����q�B;�ͧ5��e�&R���8�]�Gbx�W����Ӷ�ouy*���P��H��ō��+�m+R�*�P���U((g[|� |�/>q��.��e��N�l�ƔӞVP-4'(Ĭs<)Q+�n��7�,߰���B�Z���>�8�gaI���vP1��i��Db	m�5�d�N@�ϓF�`p�5mt�@Xa�|��O{�w���m�Qu(3�iAM2�NA��WZ�ֶd�3ϛPz���N̷�Ճ��~u=X��0�m��������N�(!���>��p��n�3f�)��j�j���[��lH��^�L�(OK��X?.c�RH=�e;
�*�Oq���0�o�e��h)�� ��둃�6����I���6��LW��2{
�ӝi��\�k 6�X�.d�B��"i)t�Yk�l��6AeK�m�j��/��'u������`���c@古�c���ٺ����>��q�O�_�dQ*qu�wYG¦�̏��˹[V�o��*��SH//bex6���4�L&�y-�Au�ɲ�txb�Ds
*�2�'Rݶ;,�sb
�b?i�/#�G^nQ��J�Lo7|��ic�6�F(u�%�2�}��M$eá��7���M��9#�u�p�~��g�M��C�ѯBЂ�n�9����f)�t@,C��E�J=DXW}9#�Kf��w��ጂ�a�]��۾�Au32n�/xً�Laj���b\V`o/AS5`|���\�/_z��4\ت�_'��0� Lԝ{���q��xgr4X�n��'�|�r����9�ֶ,=:T	�����e�t�X�({���B�
-&5�p�^�P��5�n[�]�̴O+F�ٍ8�
�\�z?"��K��~�bs�Y������)�4�7�$$��r�{Ż6����l4��4!���+�=2�C�7�f�H��3��˥�����=�s�+�{��O�b/.�@�?#��y^E��-i���>��q:������q��
�o�.�BC7�+� ��$ � =Ԩ��y�zގ=s�!��o��K'����Nzu���11,��;��ּrjpՆl�K��St:O��<H�'�QL��\�g��D`��F8�t�
���L�����L�ƙ�6�kK�W_21�,3�9��X��B������ o�nE�(o٥(�u4m��
��A��ORtN��x�B����1�T��0��x�[(�״�ǥQ�����{�#!���34�����㳾Hv�fD�n,i�m����F�*;NR�ڞ�ȿF�6=�̳}L�{����
�����E�2�RP��G��H��@'7�F��/p��6�����8�৖F�:d���G(�9o�=��v�t���̈A��▫*��UB)��ED��"r�S������"M!�qV�֘4c��[�N�W��J}c�P�������v�J��ї��f�>�I-47"X��|kA����˟�A(��M��9��RNU���s�4^��b`:�s���8]�ޮ6r����pꆛ�/3�����4�ȩ ~�H�M�ȳh 걍k�&�wfo9@Y�)�)��An�|��.�q̻�2��\�Ȏ��6l=��zQ�3��XJ�J'�����r �1���	�MU�9�ܒ~X䄥}���hw�m�`AC�5�Qx�@B��LW6��ʗB�_�:$�	Se�����XƮ>�h�->�k5��I@�s  z3C"�B�� �ɮ���0a�7=֍�Ǣ��������^�#Z`��dwm%D�I������P�3ʛ�2x��<K�� ܓp-���{���}~���[�y~����I�%K�<��`�ixU�Դ��_����.�QìDF���=�<� ���N췘���}c?�g��#�"Y]*$��le�,�(��)�D�ޙ��(=���z-V�!��H1+q�2�Ā
�cԚ�+=�A��R�`��iu�'(s)�\��d��s��O��6+���"<�Ԇ�_��	��V:ݑ��1J��;s7�9/��"c^�L��`�bH�R�����Bl�%"Z�j�a��m�J�7K�`�'Q4hRS|P��P<�[i<�\�׍��5�6;H�p��ؿ��w�n���J+'�7�����q��}c;U�X�����mZg��A?=������J7�R$��H\1��iZ�F������Is��n~}Qx�!3�6����w9����"nak3_�X�����c���x�]s�j�I*�"�vT4a\
r�ʈ��o����(�v������n�HF�ЊEg�7�7i��?�J�y5���]��\[d)��a���Lrf�`�#5���Xf��*�v+X�� �@`_^��t�iE���X��l(m�Sl��� �\��<���2�P늳���&� �n-�Z4�ϒ�t�菳l�EyN`�Udu ���kK� �:��X"CeK
�2�ͩqԓuq�P#no��l=����F�f=Z��l�
H�A�T��Q��;w�����r�Yg:�b�Mw� ��<��P��\`�T+�?S�����5}P[V����^�r%���J��0ю�Ǯ�g�ْ��E1�-��β�$�1v3g�5,�"	���T����_$��pjd�*�#�^���A�J��q"���r{��t`�r���,P��֙}�{tXO�M��r�"�����f��6���ִ\�R~���4�҄"�2�W�u��8��O|�B�1UO������&6�\H�D�(")�����_H�L���>��/�h��(�+��}�r��fپ����*C%U�ij�Y7I��������,�f�\���^�	0Tx���EV�)�+�jќ��,!���:��2v�5��&ۃK�>m~(5=)ol�zI~F!�K��� ��<m�)�֑�0;���}�2e��h�,�g7��d�q��3�*s� a;�Nv�Le�X܎�ێ�ݚ��1�$k�?%����>9�i9�~*gp��-L������->X$�Uo{�p0U! ���x5#�

����7l����E\�|�,�_�ֽҙϣ�
ā�q]x[�J����dYE�Sď��.o/�*��lU�����I��1�'K��'�9�ԗ�KU.��rvj�������V�����ӱ�iY��j���0��jh�=��w�y2�v���d�pX6MA4��q��L��O�G?����V�?]6i:�qa���V'�)��bNґt�.ײ`���-�}(꺤�s'L�����t���W�y?7���{���o��u����0MT<AL�Kn��C7���aX��)pN$��Y���j�w�M����.��b��)���J��Z� �IZ���_�yH��Hԣ{��Ś�v4�ޮ�`K�l4붻�.ɚ�_�^U�q��l�^����NQ,��{��H��C�-��F�#�7��~�������J?�@HX1���K7N2{��j)��֞YOf�z��&�S�o�@�y�ϚM7�f(��N�@��e`��N�H�4�HB`�E����XW�����;��N���4n͢ⴷ�%B�o�r��y��dD
�;�Fi~RjNue���+2�8JxVm�;�rbI*�g�;�|1|��\끵=-��r�k\bU��q�$�/�n�e�" '��'V����v�;����x���H���E�/�7lX%l�X ��o���u�,5���H���v�\@�k��2z��iP|�t)���6��x�<�ך��[*qD-�I09l�W�4��V � ړx&���5r������#d����������9�4�P[��|�܏�.�%ʙ��d�W�ˑ���C|��NlSڅQ���<�a@��(�R[[.}��-�-����G����u�]��F�a�o:��:ݢ����U_�Yh=�4�,�"U��}���[���
&I������K	M�X�Pj�\�'#f����ud	������1+V�d8�ƒ5ʜG���3�1C�$�櫬��htM&a ��@ݥ�9�-iѾF�V@a
���F�?�`|�f�҇aw�UOּ���^���H�k�p�j\2&�K��ٯ� �/�h���O�.sՈ�He6g.��O�07u���Ĳ�#�͝�0���4<F���}̤����K�Ǽ��J�����I�0�C���+�#�WiN)����؍On��H�Eg�界����t��1�8�_4o9cr3uc)��[�E`=�R����@u�9AJ��I���M��N 7�~�ǃ�s>�Av!t�����0�p�n�%BL�N-��Xr�JH�Mc����VF���|�@��5	�d^�̳��l��\�]"�~U����C@��H�Z��w�B�n�o_�1������%V����:�'�k�ٮa.O�5���`�ZO��;���B`~%�ɴ߃M�4�\_���?��̋G�Wr��e��MԚa��ǽ]�rd]��}r���%ץ�հ�n�f�A��ޗ�X�[���Cs��ޢ0�[�\����W{�Ld^\j\b��ŉN��שa�#�ɑƿz���hQT�J*��j��\R6���r��	����A:�i;�x�W����\�}Z��>)�"!��^l�%���M���{�e��Eyt��R<�+�v�����W�~Y��M��UuG��/�v99:�d�����_���%�|��"&�,���B �W��4x�5��%E�mj}�2�YI-d�%ʺ|:+ߴq� ��F̀ch�c��>>iqL� �NG��N'��E�oKl3����z�VM��˹]��J�lӾ� \��w�T��54Kܡ %ᥚ:29K8g���?�A�D�X:ʫvh����񎴹��*c����}8X1"q���G�M{�����N�-�ttAv��s!>��'��s�g�9u�ȷ��A��
 d�Go�A:|MO�v�uET����]�w�.R���-,NGW�����������(��K�Ԑ�+z2����
��l���mM� ٱQ��w�K)�'�\&+�,������� 0���v�u;������ƅ�
�Y����΃�C�S�n0��ka1cvU�Ln�q�y��}���mo��1^�Q�MFN�`�yzXt��*u/� R_(��yu��G�0����TPg��ADVX/�_T�ǫx�P�B믑�BӾn$,�7!��"B*�po*$[�-�$���]��LD����R&��u�]Ș�� ��Z��L����k\��R�;BM�F+i�.������������h�cE����<�X��ꉗ�÷9�)�]n�{z_�n=_���P�NRRU,��V�g���vz��Y�( jRo?ވn-���^.|&%*.�^/#���a�P�sC�4�*>|���j��=޾��@�p͖�߽��ݻr���"!���'�eA#A��$La$���f혀&�:?+���Uw�c������%�`���P9�Z���M1��x��8�67Sj�2��B2�J�6�AL��u���/�r��l�Ev��=J�ǀ�����׉E�*v�T�g�n�m�}�C[W��}w2KՅZQ;t�.�~�f;Nx��Hp{n�b���)�T˺]�z"����́+��m-r��GB;�y]���m����oߣq��]I��Ԡ�aqrh�N����Z/�	%M/kf�a�E�n��^�5o|%t��(Dt:�@��D�"4�hy��7�ߢ�'��'�e����a�G�q�ő�&}А%kʖ��v(�،m��s�ݻv����0y�<]㼠��}a���Z�oq��DL��g��#^uQME�Q��a$�(�Nr"��3w(���6�p�'��z	�h�����,|��R	`�p�Q��?����_���8^�����cΕ���4�Z_�:��;$<�so���d��v���4%�3GR-: ��h�k	W�ATڌ�iWo�Rs,�a�!0ѫ�0_�'q����%�dn��&���oQ��8?¬ox`dg���U��<�R�O�>]:}��qP�SZͳ�9g��n>�{�(b��>����%so(r8�A�1omP��ڠz-pM~Gv�Fyb��Üe��_5*ކ`<��n�V�ʻ���9��a��1eMl��o3 xOY�jw�)v���	�v�}}a-��P���k�7j�*-��PV��m]uYqg���H�$!��J�,��*��}!m�sƶp^4���������\V>b��ﭹ>v!yM^��Bs�p ���a�4���t�������|;��[ȴ��ȃ�m��͒�ҕ�m��b��ܰ��f��8߹�Cд���!��6�x,�y��K �b!"|����l~I:j����Wepsh�$GR���nQ�sD����9
�F�2�d��/�yq��c�T�,��m7���_l|1�-!��Z���$mL�l����ivB��Z�(�/���e>�{*7k��ۼ/#��9cr���;d�JA����1ֽ�q��+Б�AS�l�\��ϟ�	���ʸ n�S�{;`��)MA�e�䭣T+���n���_\�7�8������Ms&*P�oUU�91)�Iz�0��F]�sJz��4�=�ڱ��x��,:c���L6�`6w��$��o(�Zx{�9���T���dB��J�|eV�$��sk���c��Pg�E��a���m�!���������o9�aV}�;}��I�.��(�o�f���|6��%'����ٖ���Ѐ������c��?����:@�v99`&��.5�$r��P%"ݜ^���׳��^��3z<�oaD�g��I�x�!Rމ��&d�P���^�挥zE��۝��2�s ���<�~� �#����
a�GCU��)L�gx�Jm�r����|��5��S�di^d���_�+Ѿ���ؑ�%��`A[�l�M�cN�tG�bq'OC{���Oݥ����R����#���	�WB@�WЃC�,�5�@���W����&l���>A|:3�d��ծT%�<d��T��l���E�]��44��`���@+[,�l�̡k-W^��v����y�T�`7oSO�Sfk�aY�eY�k���e�.V'�߄h����TJ?~��1�%��ȅiqe��5�!��h-�8B?�E
�cL�� ����O'r)���&��[�^T�{�?���Y�u7������.��&�����9;?����N1g3.Yԩ�%5�Cƚ�*�P[6-z(R��]zp��9� ��@/sN��3�K�t!�03T,��>e#�ɳ%^�0��V�s�yƴ��+��70��Gt=�˻%ZT�	���Q �@K�H㊗�X7Av�{F	[� ,�{o*���ˊ�;dV���J��b�V�a���1�=U�د��8i�er8 ��el�L6�:�ID�z���2/(AV����?j���dx��Փ鎚g��#d4�u�������Rs)�aU,��� ���LB�kr�~��:� $�����{kP��MDyr5*"'���3bR\8e)MYR2<�V2��ע��Fe�G���B��Ե
��?�BL7T������~N�$��(�!������x�K��X�� ���>�҈찵f�&��m�Y�Pd^�aW�O�W�Jؙj}���-^(�d�xF��q�9K�a����)����o���ʶ�ƒN��9۝?�52�˺��uf��NI_�x��g?P�n���Ή�3쎔��OSvxZ����?&w�"=�lR�4��|4ȩ蒧%,r�M�i��Xv�A%ۿ��V�ͧ��Xv
�x�#�ȭ:�q��-��B,�Tì������w�~���������2�=Jb�"t�R�%D6�������a����0�j5��)yL�	���iS�eܜޫ�\?�̳8I�ߦ��b?��s�^�o�s��;�ؽT4ˮwN��E_.�\/s��r���r���Mhr�smYz��w�4pX`Wu��PHĂkNү,�]@
;�#�a?w���j ��=���S.�J��z������?��X#p�?��B�g*���/چ�zWc�qF�q��o֏��8:��,�~l2���tS�1���J�ؓ]5���ն4\Ҩ���o� ���;y�`���@��)ˈH�W��]����Ӂ�)����b�zg>�>�q�<�$�v6�3�Td~��M5d@bu�Ƹ�kIg�}�ii 9|��C�8�������+�?=@���v�S��Q���H��K�hʣe�j�l�N��h��s��=�����pڨ��x����[�ώ#hbMZ]�NN�����XI'=|,_.vq�EK��R
Lc�k���{�u^}��I�0@ذ��H`�1	(�x�ֵ�nz�3�S�i���=�7�>
���2r���E<Z܏We	4�%���o߁��Y5�B$���*D���{�J#���R���)�6}w)v�u�e��l�j������˓�Ӂ�J���uiG�(�������RrȖ��P�਑��T9J@}�=��j�BO��k��i�����\k��N��u�F�[�>���^�8g������w:o�u��`�h/^q�ɹ��Fi)�M�=X�z�8��Α�ɳ�F�,�a��.
�����Ԫ��̝,ti���")^S����]��:0���ը�bj��zaO۸ދ�[��C1W�ɉ��Y�-�.����.���b�1`�H,��=
�zd܁]� �S��^�ր�� h�����8
�>K�N'aY$�W�"� �a�����.SGH�r�.}��c��2�ɗ�;��f�xC��B���|��5f��6t�1"�
~x������i����ސ٩�������ܨ�����ʓK;J�2���M�tÄU-2��aK�D�\���/��2[�\	t3�l�0/ζ�c���I�R�w��\MxR�ߚ�[��	f��=ו��+p滐�S��H���+­���2m��C�0çXf��G��I��=K#F�)���$nz1����aCͫe�$���|���H����� ��E�Y��|���Pg��^5��P��y\��y�X��51�6kp�mj见�����LN�:��d
��hn��*��iu"�J(�Xƻ�NU:��ϧ��rW�e�얒#\�Ƨ�"��&�t-aF	�����Fy��F����T��D7E��cLzσ��s�4�J��T�r���U��'�$������^5�l[���x�N�u����Zfz̑�Ƥ-!��<�����*t?73X������Q�t�yv�y^��CZ�)�� $�+�]6P�cT�F��Ѵ��D,��>�>���h����~+"X}S��<�M��J����v��x���5���Z��	~ l�(<�}��"u�,�q���:8���U��ˠm�����4��ZZ~q�r���|گș݉��U�)�i%蓫��PDq�Ȩ5F7���K�Y���u�Ezk굵�� ��MwxzP�'�5ʆ�@��aE~2g=z-ԓ� �.����֎��L��}T�<)�G���9J��}.8Yڏ2��d��_k� i��[(»�s��w���#
򸑝�M!����ƆA��Țr_�z�cD-��%���`b�:(E�HJ�6sD�\��3h�B����=\��8�_)���5�L�y|��wߤ���4�q��1u�0�������-����g�D<��[�VY�A��T�{�>��я�߼�ZD�i����u�l*�j�a�I��h�T�O5p�5	��q�
v��w~�'�MN�0�@�U��	W�ql8���k�:�t�
��N�꘠�$�"mat���Ř9��
����;ft�;aF0ҽ����U�^�â����r.!v�CG�@Ӭ}"�v�.��d��®���yn�0�i��j�sɪ���,n��>����ZY;I+Y\ާmZd3���ip����*~��v׺h�OP�RW�(x
9ئ�S�y9������Ş��<r����H�����K�i��r�ѿ֤����� ����e�����*�`v�t�����'� 0�rcP��c
�%��{���]T���^����������1"ҳZ�o=ܦ��F��A��}'[��V�h,.�$րO�6M��?��j��B�lEE�f1y��qza��vڐ�����R1����\���E�ߤ�>��e����P�/LC�{�H� ��R�-	�{8���<����D]q܏�$zz?J���X5}�J�����T�;�(�T4R�I��0�F[-?����N���o��)5��!�Q����8n�&Q����K��I��5�f�D��V�e�Q�� �k�Ir��3od`�	
T@�n��U=�zE��O��迤�8���B�Z[L�����12C�4y�G���^�� �1�w�b�v�h�W�k���/�康[8 Լ�Oĕ��KW����"��?^MqF��~TB".�g,V�t��R�j�}�dLR�s.&���#�X�PY��?6o�;��� b�z˾a���8�_4���}�G^�U^�#�G�n��Ega���BQ���~z)++ZtGN^��Y2���=}~*�	œƤ�"�H��� a���T��r��v�
;55��Q΀�f��{b�&�t�7�����88ı43Z���UH##��!C(R0�� 멫z,�3��t���x��W=_�n��0��+ĥ'�	������ɲ���*����Y�oZf�����[��8"��[Ok�*.�UC�����W�Do�<r�Ǘ������uY7H�|����a�P#�Ϩ����*����*���b@17�GT1�����������-{��D4��$f��\l��\fhբ�A�|f=X��XTǵ�]�;�@8�|�[*qZ�˲2��5��D-ˍ�ȌC�<v���ZT�$.9ȇc+�-[��g�C-`]N	��U ����#M��I�EZ��q����Ѝ��ݘ�n8�(Nߥ���H�$�s����" �1L^���x�ἇ"��l���iܜ�
l�פ�����E�<����Ѕ" �x~����.,�M����)m���H�é�����@������C#�]��[K�;��[���1B��>P �}]�bV'����E<�G���ˇ�a�Y/���X��m8G�Nt�K�
�"ٛ�{��<�ԓhb鞾����g,
����W�/��40T:��YH�۴����GQ8���x�񀈹�}GS��G0�R��NF�T��C�݆On�Xž����#?JQ<>&��)ü�H`4�����y���	���|�N��1� ��9��
���j�6��)�<7|;�(}X�s�pʞ� .�cn���Ǆ�m[�W4؁"�.K�v���\�y=���(�U�OL���Y�7�ʐ=��3ۼk�.�V�V���q���s�dO�p�gL2VR���R
��ԈX��;E�3챴�v!���u	�׼��ȟ��+��I}w4��~���7{��y�\6��Is�5�IPvv����G�|T",����[���)0�������CI5�!|���qTkJ�L03��]�������)�-eg�˷����o�O<�v$��P��:���,��H�n�6T��ͻ�xp�u�	�j��/�}LX�߰d/��Fz��]P�)=Lus�e�",�i3z�������#��%�`Vݮ�E}=ec��������{yW��, Au���������n �#�U�A���^�?�oӳ_��K�3�)L��!`9/
h,�bʬ�� 6P=�z����a<8� ��u!��$	���w�Ou���:�!TŸϜ��Q��gF��s��a
�(3��͗G�X*����;�vL��<�3���߱Uy��^��R'xOH�3^�=���k�
LޣM]�����Ԝ8��QZ=�v@��_���;���/e( 6����fvߠ���Z��L���&7�:�B�rQ���fԂѱ\O 1�0��9�欞ʼ��YV��j���P�'���>���^]�D[	�`7�/JX���xnC�`�?�zzg^����hBZ��v�8�*yS-O*C8|WR��Z޻y0{�^��3�� ��q��e?Ч��m0���"�o�zK��IUk�4�|:-���(B@W�f}��I��w@��\?%����E�/��Y���^l� �|��]r���JS6f�����4��������x���ets
-o�?���M�+����J����� ��\c�ƈr�ߑ�"F�#�t&��pٴ����w�������Ù�HPFX7�|7��j��7�=o*�$�뙯A�q�>C�2�~ψ��l�2�;�^nc,��v���d��&�i�XC@�5�<�,Q��X��2�8}"��y�!Q�	Т���5�h�S�d�����Ѣ�Q���IQ ��Z��:bQ�y��Ҵm�`�$����:;0~��a/�F� .�f��h�8�d�X6(d_@��hK%���:�.c�� �Г|!�C<N�ɚR�Ots�c�l�1Y�W�ӺS�p:�B�L~_�-d�\�GK��o���[��� ���,v#�^��w�A!ϻAYv�Z��ݚD�A_[�����s�ңdX)���$�[��~Y��Uǈ�5�7=�g��V��F	��g�)��c9p����ǧ��|R�%�{oR+X��`C`ڥo��V����.P���8^��N�)�N�#�� #qk���o��0�sٹ�/���jk�G
6h����ײJ4��I������xﻳ�Rj5ۓ8B�ή	F3�>"���\j������T�Y =�/����wi�I�T;�\uZ�a�?ң�8\1_3f���[u/~��̻j{��z|L߃����Y�j�mR?�}�iQuC	A�a�L��Î�<�,�e��	!0�'�nw7���+�� [!�7b��7��ٔ�<<���䌞kY^�x���~P�GG^[Y9;�{�n�����ѢU�\$������фd�!�U.+p��p���\���H�X����y���a.�O��?�P����X+���P�8��О�4 ��)����a�8���S�Rs��A�P����?�N:�P��$!�%�e �wo���"p���i�����,U�y#K'W�H�(窱�9�@��I利���@��mXE�eX�a��pY]zh@벼�@M3��K�R�$������}B��x�0p���lS�����[&"�� �	�kS#c�*�x�Zw/�+�!�R�R�S�.�F8�����eG����I���mK;�^�������:�&ŵ:kX�_s�.���JPǱ�x�0q�PI���HrĖ%��L��V�눆�Sy~^z�~n³"Bp-$bI5��鷄���y�(� �i�J�^$�C��|hS�%�-��7�u�%���&�����sư)$8?G��=������b,����0�Li󘴿\۷7!�풥��ؚ;�~v��Q5O_B'˳e�y'w�K�ܱ�+����Qbrz��L�֙��H��w�O%1+BW|i�?��$���s/�o��?z�����ȗp=V6�LDU�z��r�"KF�=��L���D���35��� �5�1!"y�߹ݬ��O�����0���3��{�(�����k��Q*8���
Ffd��a&Ke�����eΎwѧ(��C_v��*�6Us�UV�:*[U�n=���#Zk�8��F��ґ��GA�u�p}�����Tk��UW�d��L���߮�H�]YV����H$�W�nE��T��0c����D���5ǲ\Xf.Pn�R�Q}��ϣ��Bt�j�Vs��K�K��>����7�8M�s*�2hX�B�;��{�Ĝx�'o�D�9.G�䆀|]�|�i���'��f�yU�e+q]��!��/���x_p�kJPm�%S��=�7�?�>�}m��g���8*.~�G�=:�xL���fJ4���^���(*�C�C<�R�����|�����;t3&d���Z�+'ɋ�52��(dj�w8�����^C��nj�a�C{�b�4�+�X&�63���d8w��6z#upȖ��[�=�.�)�����#�@n���|�����Y����i��/x��i`���Fjی���aG���u�o�*���B��Q���B'�!Ds��K�q�"z����E����=iS	��b��$�i�e�6�����C�_2f�!�����+��M���	�14Q��6u���gQ���� ��&��=����Y">�M"����՞����������N#\�J�f�W0�Uk؊� �Mc4�F�q�5���!����"�-)�/Q�4R2��BȵaJR����2�_��,��ڋ눖�x��y�`/�w����8>/�

�<r���&�k��Ɲz�Y��s��֚x��j&��L���:�3�nt��dW�/��F���Ge�+F&�C��R�S�	 �������<��7~���%򗤻t&�L�� �¾�o�2Gɀ�{X�,CV -��<��y�p������[*�
:�?	�5��?�z��L{s�٩�7b*ŜK@��ʫ���'I8ZD�=p�މr�/�����ꅫp�Cv��;����.kg�7���M` ��t�'��w�|ܷJ�WE�E�7'} y�p"H-���.��$S�T�L��t�Q�c����Đ��g�`\ww��) ��@��2�J����[�W��\ՙt�!��d��/a}�����b��l 㚄 ��P�P��}{���-�qRх�RՂuR�J����!C�q�:7Q��M�B-F��-%#�r4��������B\P�z������n&yLwĥ?^&�r,xy�;#�]�	\��I�b��
�e��&��Ot�&�+8� ���y�F@"�<,f�6m�M�oxP)����҄c$�ۅɁ�L :�Z�!������s�{�T����O�7��aVo�uo��7N˕N���{�������e�o��<��>	�W��M"T���o��Z�g����f��C�>ni_M%�H���tyd��������2bO��zvA
VG�g��}�~�{8kVX��.w�)�(Z�Ҙ��eN�W~��%��F���-�t�!��?�	0�@/&[�"�Ӽ���udi��\T��v�r���Lcͅy�hݘ7Ѧ� `|�Ǿ)dI$��C�R���$AI�W'3�Us>��z(��ޣɉ�g��}XZ�ji&�a�.�sK���xg��K�*.�i��4�\��y�m�M�,V�6.:�Ǘ�T��`���;�����ywI��!PL�^��⍥٬�jۧ�ێ�
?��ma���siI7%:�}(��=���Y�+�g:���b��5�^�kP:`q�}F���k|�(�S�B��ZV?���� '�B�f*y���>
i�� ��rPf���[� �6�$x�̢�W��'�l{M�[����[O�'�{ ��v������O��*4i+A�|��I���+��8&MJ���G�{�||P���b�[�R�3�Qat$��bl��WV���)}>=��e ��7a=�[`�a�kވ�W?�N���뼟D�q�|a)���eY�dq�%Q�$�ϫ���|�8=���ŅU�/jQ
Ye����ͫ\��
${8�Lq�#UxsǍp&��;�h?��AC�Z@���`�}�:�l&����7�<�����3Z��<XP�0��Z��{u�����Ť9�W�y�]F=	�"	��_�~Z|>��"������� �kYD�C�苶�I6
�I�2�N҅�q^�c�������~�����0e����2��h@��Z�*X<
+�yl��^���vH�}D4�$8�r��7R��M��&��3d�N�<��Y����8 ��H��ؿ͊��q��o�Mb{w�X|⫩���~�����Z(�6��?U�s��Nt6\�8E�%La�\w�O��)(8�t�fi!A	ZۛAߛɻ��E��,�{'�g��]�@�f��|����v����!Q��[�[ӋnFA�U�jes.7�����3� ���k;_�@ˁ��z_Rǝl��ޙ �.�.��'w�U�M ��Si�t�Y�E��C�O���}��w��4�%�>$/.�+�O�l��b=��l�� @od�T_܌=��ͿG٤�~ĩ�AzZ��лQD��#B� ���~�*=Z�)�-l�*�+f$<��b��jN\�Eяޮ��yf�ͷ��@2��G��)���tQ��������`��!2����إ���A?$����L �a3)w�f5��(�qx���#�d��~�-&�iN������=�xa�E���&��7��/�h��V*�V{�(W�Q�b�'�=؎ˮQm�V/����nO���r��{�~�,r�����P�<�Ѱ�Y _�q��D"9�'� ��K���t�{��X�Qڥp�8�5����	?�!����bƭ+j|��X�:���v֎ro�c�R�ο�����j�S΀.Y��57w�_JwC`��3����O?�-��O��$"B�lt�o��e�	(!�39���*��	Qj�V#X�3��&����bv^���Y��@�
�u�����w������l��?$��{�� H��_���Z
	���v�%c���	�d��r�o�{x��f��`	/O��U�p�2H3��w���ص��Yu8���6ڮb�5}y|��D0�����J��ͤ�ʔ����2'�Ե�`M&'����̀ԅ蒩�ۇ��w�;7�tGi�z6<>�������r�Ԑ2}��h(q�|�̵�1Hu6�ݝCΕ����%#$mxB;E�p��鎀 @�D���n��C��<nx�	EE"k��cD�&�lkUd[H�I=s�S�1o[d��xZ�]w�����X�hDK�p$Ը��6���Բ��;CM�"kc=2��h���K��z�Lұu�EFT�j.�A�3�J`e�1�ى{�����B�t��;XlGp32E��Δ�ƶ�n[����� �yE%"T�4;��;�(��H��z��W��EW�;�t5@����p:�rS�>�:Z_<ఌ��`�vt�u�w!w�M�p�E3ܕ�ν'���k�!�ʬo<o|>Ke�bk���O���s.��B�i�&��0Xٛ�o�C�S`��l n=^��,�"��0���S��:��+��{��s���b>̷~<]���vS`�ڍ��,�Ǧ7FG���o��w�Q%�[ �x'��=��x˔����]�'�,�b�fD����%�ZgM�k9��<������F䁂�S7#�ʩQ�ݻU��`���g��a�#��k��I���@`T���a+��l�q��B��w�|�i+)`��N�K5�ݓ�-���������Q�e��tϙ_����c�˞V��@��^Ip������3�jFkz5
�˰!�|n�gz	h˜���nRG)q�k�s�GXѣ�ݦ��{��ѹ	�S���3�d��/ ����
`�4w�;�	<vi�s4�{�.J��:ko��tj�}j0�9�n�.r�~"g1ޓ�����̳2*Lh�|^J�g�+�^�kQq��l-���ϒz͜�p���)��?LX���As���%[�b�sHi����A����j�t�K���e	M��΄�[�7>���:�g���/��IB
dDĥ�)�?dܼ����j��Sӽ�����:F[�r����}s���%�
~o�܁þ��n��a��L���+c;L��ޛ	p\��Ja	:sFɪr+(m��>�s�̓F-��.�����*��E;��V�'�(�oR6*ؒEa�C<*�q�������E�4�/.�{;���,b�3u�r$��';.����_M��`���Q>Ip��N��#I+*Z��,6}��.$u�,L9�qh��C���$2}<��.�),��I�ֵN-��{Ӳ�V?��������H�&5@|x̱	#M�kݟ�MQ]�&H|o�1��qwp�(�K�*Sj^�w�0K@G� &����n��J��`%X�C��|\�2=�#ί�СXV��Oo��Nh6��� 	+/iY;HE������v��E����S���.�t�6��w�J�O_�e��|b�i۲��0&��}2E7�Y2#0���D��0:LUSh�F^���R��ؕh8Y@�̎�Q�!�ٴ�L�'�k��T*b.�s����3�t��5�qR �⏾	۠��EF:s�
n�"ƷaR9�Kݕ��vp�U|���'B������-5�W�����Gʲ�2�u�o�SEͣ�>;�_!���C�C�E'�����w�A~�ү�A:�����/����3B[gʇ����{�i��^�wA��������M��oL6�L�!���w���b13g$]ɐtl�����3s�wغ�$oO��ꈣ����Z����&2�S��� �(�����R^Q^�~��]�r�KJ� �*�.�a�
��L_�潬�(���I��"X�[��K_�Ԩ��@Pu�L�\$��F�J������!�+;��u�A�1�i:&Hc���8�=:��I���MG�ly-GY�ﴛ�G���,������� �03��NƝ�Җ�ե:��bi1K��J2>%A��R�餤:�{��T��o!�����|�gy�si�����/�PK��j��x�%s8M�B3�R��e�o���uDm��X��:9�۽~)Q�Gyz�U;d=#��	[[{��H��Q&Oc2���_J����|3B1?m�$'���t^���ۚ�<�]� ����7���P�@��TWiM��j�"��;/���VR?�2p׭�B[?ЛzO��T�]ɿ
�V�����n�Ġ���/��c�:y���uG�S*`7�k���yCݱ�oH�ϱuB!�����$���;G�i�)������՝ȎJ/_�(�h�U뵄�E�W!��PȾ��a�
j�����ݷ$v���9lu+��sK#7b��R$f5yh��D���4������U����ox��T1���@L�/)h�g�e�e.��v�+����N�f����w����p���g!�}i}XcB|wbC�4�3�����|Nަ�b��}z0� 6~.8�n����Z^f4���3�U3�=�]��$ZvMB��9�N�0��nz�e��\$�z�-@_��Y6׭�BVPh����Bk�����u�����Y�p��}�+l��.U�j"�y��c���ۃp�;6��궱�(��%�4�#�fS**e�+��L;���$A�M*\1�K_(����?9�Ç�'�;T�\�;i�*�����}�>neq\ik�	��������'(ODs�T:��71&Q��4aV_C�&����2��6-�]�p\�{��/�)�;Zcsu�V���?[{s��X�+2�So-�2���h}O'�?��M���~1Kf������V�P�.S��u�ƵO%��#���N���~������qZ���E����%
q7|;@@�L��f #}���#H;���H�� ��B5���#N�+���Bc��(�se�ġ~�T^�7��h-��%;z�+�U>n�'J�B�Wﶙfv+��(L巆m2F\��n��ׄ������]8�hN(`�����f�;B�;����'o����=2���U��uO�G��*���zfUݕL���G���^ �J�3�^��]�n�^닍��1�,���dt/�d�0�Q8�q�ޟ`#?#��6�f�����$yS�F���va��o�fy�&�,XG�/&$dƞ,n�qO/'��V|���8S�YH#����_����
(�\�к�ߍ���v~^�L�I���hV��&uC���UgR�8�%Q�dM2O����%$�IKM����*M��&�s���i��*}��-����w}E��:b��w@,��^�#�l���=D��1��J��aG� 9.��y�����Av�Ɔý��N�I��?�I*n��O*�ګ�;U��UUk����ܞ��0j�"Rj[/����\Ȼ�o>ٴ?�Å�A�AnoOfº%�i�����Q��J���ߠ����'6�8��[ ���� ���j�E����Y�0�����V�㷾�#���
M���T��D��#5��D�e�)�˝�Ȱ�t�0�{���G)��A�,򻊬��!,��Z��� o3\��C>�o�R�JMg����Ⱦ����;븺��#�W�c�?]v�����p�~J���e7W���ZDw?�3S���: 7'^�i�T��D��>ޥ �F�|`Y����9�Kh�Ρ����ƀ��46�LK`�.��&������=�%/�Cͥ��3�8Vr� �&8�~�vD)|��d���b�G,�:�Z�F�V3��L��@)�׬�I@K7�X>m�i�1E*�L�7��f8��ޚ������b5zPi��Q����IEM7���Zb� J�E�íI�<�Tu��Ow��a�[�,�}��n�_������ڋ�ML��+o.4JnmY��8�J�_[�8������!o�[�0�O�Q�g��Ȕ���J$齁��>Og�y��K>�����@�/XzY�81������K(?;�n>�w/���r�t+=�^�|~�^:����=� ���d�)A YHe�\@��P���)�B���t�ԑ���+��G�{K�ҕ!Pɉ�C��;�r��&_U=V.	�}�倏
�ᙁ�z���.�s�BF�����t1��Mǲ�	;�������.*�l���{ӧ<R�@�6
�h����+�C�n�����j��l�+�#7�������C����|���ޫI�(%�� ٭�`�M�zr��}���5;V�j�ˉݴ�֟�x��p�n����j��$�%8!{�����6�;���jK�����}Ua�bQ�0�Y\����RY�h'����3�I�$��^V�_3�l��r����m,���������#)}/Og�0�O?s3َ�2��ѩ�VWi��c�)��f/u4�˟�f�),�x�sL6����/;{���\>��Ӟ,����Â|
�z�5r�ҵͩ���)�����4͆�&Ѵ��/�DH"SZ�;+���u>��{�z/���c/���R#���9DtO�d���#�.�9u;����k��"�EW�O�J������|$�V��X���\����ře���ީ�3d�C�Z���`tߴ'�)�>9�/i��h#�����:�+��I^��J��R�����^7. ^�{�U�w��������(d��Ѳ�v$��MNC�F��I��=2|���N�O�,=5B����ǃd�fk���Ɲt���,6�<��&�+��`��w39�	3��dݯ�c�_�x�e�p�6H�bE�Ct�IU��{;)e���� oz&����h�WK�k��=�q�|PovMa�]:�8pn�.,��4�����9�������-�>���k�'�s���b�+�*;?�#K'Zm|~օ7_fZZ4�e�;2��E�ep'���z�lL����$5�D
jk!9�m�֦���|:�SF7cI�S�%t���S`�y���Ѿ��p��yLĎ��R��of�~���EL�o�y�Y[0��^Y2�g�Of�9�"��ec���O�]�caV_�v��	����l��	@f)#��_Y�MLh�D�����煋��@:qV��2']�1V���`�y9��K�o�Ojz�(u��r�J����I�E�C�`��Q�7y�ت�I8Oh��f+!^IO#lt(� �� ~.��CMe�w,,�������R�-�|�_x�x�¨a��&o�W��郮a�k*�,F ��z�^}�A��i�g��ʾr��I��H+ބ�lڡ�+�߆iku_���ټ���y���B�{�L2�	�p�3O��/�[���S1Q+��Ң\l���6�[�R�t꒨ �%%X�һ;����
A�0I�"�#�-��6e%�k������ٝJL���r�V�
�>���Mٯğ�^�gW�s��<�-�&�xL	N#���t��d>���D��1ja�o1/�_`;U0�L�S1�A��*i�.�%�I�� *
�����/���G�Y�C�0�����E�<�dsA��ܔ����<]����?���q��|0cy���
��;Eh���LSj����/�9AЗ*�xm3��H��y ��_��[����ZT8��G�V+n��q���]�����-{��巬�l�~�Q&���?��'km���1��	�p����Y�z�LVQuEAH��a��{��A��M&�2�ldk���Ü�Dk4���������8�NE���Z�����;�5 �fE�_OvQ��nN�t�mb�?�.[��(���Ϊı�/jY�a,���V��L)zX�U$R�H����r4��M4u�<¯E �l3���f�+�渃?��z��"8dG^���e?�I��o�������z̝�d#U�A��v:��'����L��~���g�!����؎�}c�΃�u�̜fB����)�a�Ə_Tl��OڞC�od�21�#�,i�O)&��VG�2~��<"�N0���W��ft2�4���U�ǃ� �_ʴ6��96�[2��M�\A�}2Z�ƭ���L��}i�
?J�Q�B�!���]v~g[ߎu�q�3�7z��@��PƛU�#�M:��ߐ���@�ZRL�\1G1A".Q��� ���hN�b�i깕n�Xy�]A�|�/t�L�4����e���S�89�i?C�mw�������b�sj�����{��Z���"�<)��[/���Y��&�y�g0��AF��*�k�S\[z��4�Hh��O�ڇcB�؃G=�����M�;[Έ}7�`h���,��pb���Qr�˰���"*��~T|��X��j�N���[:�J�ǂ�Kp֐�s)ظ�	��r��(>R������쎷�L/�����s�r�v�x�T����YvrX�J�[��++`����S��TR�̽�j9ͬ�o'��	�>X�:���վɈ(�̍O��=��w�=�����"!�~��|��?�@��X��*�q3�h*�<�*��[t~Nv�������x"�x:ŭ��b�]�?ۦ��L�{�f��R��E��I����G��7n���5`L�N)�,b��v ��D��6�����q�ڜz]�5�-�hu��>�����|��O��T�%+����UiJ�w<��9�j�Y�Ow�E�_���Y��Q�??Q�^�ʾ�s�7� "��?�eV�R書��a�Nt��.��t������QoZ����0�`^`��t�e�I`"�J�Iʭ���W8
`�+,�폁�E�b��-y2��&]�V@���-\*,^� �N��8���t{"o�W�bŵ�y9t�?���Be�b�D(�Kڎ1 N�;bJ�QD	���]��7Ł"��{t���_�r��BI��@M���ӷ�����v�
�Mָ�(C�GѲU�l���y�fb��4���5�]/)W��$��9���
VK�	M�����mL�AŮo�\ǐjr��d���70u�$�1c���^�%
�[�H)m��rhgY���K��
��8��տ	����b%�ȁd�-YbC�u�R�g�t5:Ohs�B�S�"��\/.+b�S�{�i. +!%kW3X�ׇ���M�hO� p�.3uZ���v��K��&��L�G>�<L�T��T=�n���-��ˌ��J	�&�]��6�����a�C;�Z�����7��A��P�ؿ^����Փ#Q����gq��%���\�[��S�QgV����	�5za�t�v��#(�s�p�b�O��)Z�o�7Ea���~&K2�s���ok[??{,󉯧&�'	(�pvb_"��ο��3%h�k���4hnv��8�|�4�r��m����*<�#wP?�<躴���`q����t����c�ر�h67w��+��Ϧ�$˲�f� 1�i��QX#�\��H�Ft�2�S<l�m�e*�T0R�� (����=X��8b����₄e�eZjF�/���Z�Z��vdMS�*�t�U.d-ʆt�#�mӓ}���)��=�xׅ'>n/�������ũ�,�0|�h#��A6�0;κC苫��T����@7�x+���or_�k���]LB9����䞔�ꭖ��*AȘ�7��~�'r'�|����(\���X���Kc��S����`d�"Q|�����i�_'A�=���@������h�>5���9�H�`&+Y���/�&/o�t�'�����[�"`ɐ���W���k�Nb��=��.T�;�6S�� H���M�zc�.�$����e�DD���l$��?$H�ܵ5\��`��1��D��8?�z�iSm��h"��W9��_�p��z7��� �4Ѽe��c�XḰ���0��\�髳V;�̐�qn����S?-:�H�V�A�p�9{)_�_���.�U_a��@�X�ZeOM���X&������{���&3=��ۋ���EO/1	�yl���P�O 3t��:��%��j�=�7��l.N��u���o���@�����ܷT��iJpg�nRMA(���YL ��^Q��Ĝl2u�:4�!�#4[")T�q-��~�]t-#r~w��D�t��#�@�A�e>|\t�3l8�4����)6���!ٞ�':�2�5�����_GH����KE/�۞���lWE��A���st�'@�U~w��l�ιTT�@�)��A���k憁@<����D�����4�$�+�Ai�@�D������X��=�,@�O9����IӮ�r6:�@7����?�w�R���t DY��ػ|�X���)EQ�:�1��\�����R�e|֨�a��j���P�گ���D���nÓ�Պa�KV�l��͉P�}���$���e�r�w.����]�k��	<hZ$_��N�Y�H�U*R[<���8� ��h�׊wiP���#u��Sz-&t�,�����b"�}�A�k���q�y�s�.���kȗ��uDr[�s��f^B��Y�~I�W#�	E���� W�pD��r��^�#�8�s���	4��y���?��$��(c�H��)a?�Y�m�\Q|��D���C���x�k(�Q�bW�Q4�]�K �=��W&	����"Mo�w�x��k��Hm��@����B��?�E�fs8���>��D���Y�Ly�.��8�%*���+d�0�&�W�������҈&�1d����&U�`�W�ֳC9��>W�M�)����m��'�n_�ei�h��ȸ]�G���*��olZf��&��7�p���Kn�Q�!"�gّ��*zǿM,��D>p�P!�[�Ԙ3�o�Y�YX��Ι������#��6����\�$_d�0B$"�}~Q(�2&�����
�m��c�L�\tu�%)h8�c=f�p01;M�֍?Fx]q�:<�zNL�����Uh]�zm��<�D�7�zte�X��dX=)��"��%5��b5��I�d���VB���Sڃ�#�D�
�=`	��K��{I��	�`L�+�%��,��d����G/��}���d ���˻��rv��g�,N��*�.8�lS���'J�T�Z������c:9.�5t���������tm���=�g�m2*�Z��>��Jh��a\PPϙ"X;��J���l^Z���r�CJN*�K'2��ex�K�����B��(��֭�l�s�o?|��ÎhB�ߋ��Ys$�"u���PTC�d$�ư*5/�hX�1b�
*�{�w-x�i5hHP�AH71ٺ�,�� �#1=���.��p\J��1Jnι�q��ʪ07���h�(MJ��Aϟ�j����k�D����pn�m��o��l �g�|�=���ئ%�W�qCʖ�z���̫��S�ñ����t���j�T��4�R|�R�Vc�x����p2o� ��p�'Y����Ƕ��v��x��!�mo'�ح����{��Q��r�	H���#���.Wl}l��t��7
xV��.��.�;iVO��sd<�%,���rK1�@�y��#J��n�4�x{��"��A�g<�>b�p��k�� �C,ʙ}�$f힊_rk��P��	q�-��pj��a���8�zfy��� �^$5�����&�7�0���EK��T:�,�#u|Q"I�K}�f���Y�J��q.볜�(+��X���cH���*�O�"놲�'xmlC*td�<�;��!��S�^���L�7{3m��OE7��B��Ϲ�Ҝ��
��
�֝��'���h�:f����En�@
����iY]�۲/2鉍���"
��'�%�m{�;=H2�X f.?}��2sp�A긽Ϸ����G=��D��[v(��9?��n�L������Ix骼�Q٧���u@��Q�_�1k�q��mۘiF+�a�]E��V��іު�+K�!}�@8qy�GV�H8̥m�����j�@��w�/(��=��JU�-S�*��=��n�i/7[��[�DW)� `�.=k�1<W�<F�J�wn��������m#O`G�ms���N(\�bra��,@�/ƽ����ל���O�G���]pH<�L/��]��I�l�3�j
���d�A��3��`?�%~�a'�,�De]�%8d(�e%Riu$!�r���<WF�D@�qL�Mpo"f�mf @�eQ��p@�-v8�\	c�l�	7ƥ5w���KEAt���F��}fauG�,�b�?�C����`&�vx�sr�5B���Mo�6��U���S��9E_�C��:	ۇ�{7g�/+������ ;4Ss�KQ-�:�=C�&ʁ�y�+�rɞê����M��g9P���<V"�?��Q}ָ��ذRg���۵��x�zm�D�'1��\��e��b+s�d���(����ʁň�����iK�鸹*;��I�FJ� M8b�
�aO��ti��Ј�Ab�����Q@�`X6t��t�a�۟��������C�NCҗGZ8_�����.�4���u�? ,^�r��B���U�b8����׮6$X�2�,'M��M��|� $�r��ϒ�9��5į9���o��(A��m�ؒ��i���|�}O�o�M���e������~���5����;y��rhI��E�<"�?m�J�`'�&PWu����#��!mN-�}i.�o��[N�[��r'<i�C����x�-�xbs�⟰b([����Oz)O/J�k��v3�[����+W�rq�9�h�t��H��c2/�����mS���0X�BXz@���U.��d��3�!�>��$A�+v���ߥ�Ź&��Ti�;fI��.��)���pkM �q),�Co��b�t�a�[��X�v!�KO�f4�� ��E���4ȃ���렡7�b*� �%w��a� [�F�-˚�>Y�b���Gj��
\
z�a˕�0����� i�|���"�P����Gn+<�	�m�X`1��Jg*Ֆ޾W�PZGr�dk�Q9}O����,O5(�ڙv�L����15��4�ܷ�0ΡP�Gm>hs�9 ��F� �+s�w�Y�9�s	o�t��+�LO�E֊�RVb�u�6�Z/���*���тI�2� [�>����v�
Q��%��} s���&�,^K����М=>���wlI�w[��e]�%c��w��'�	�7�j[�M_Fҹ���,Y��#�:���D4G��$�?�����)�T	�r��A�*D���?B;#98�)�j�}�����<�Kcӷ��حL�Y���Ձ6U\��t�֊Q�����%�m�-�(nn�$C�����{�o�9s�N��Ȩa���Ӥo�OO���D %�'�{˙��&b�X�0~��`|���C�Ѩ�{����^K�l�NN��Gp�e�a�bö�D�t�#�3uy�F�S뾚��.s�y���fC���Yn8�kөr�U�<���clyNw�bG�x!��jϡ�0��Y��/�G�S?^��Rz[4��5t��6�n���z �Sy�A X��CX�N�������<�"�)[N綠#Ǟ�nd,^o��Ԋ�f�5�,4ؤw&�N�k x�-S�H�x����=c�էp�x C����Ƅ��-塕�ᰆ�u�H��y�;� ��.)�ֿ@�:T���yA��J��%�%��6F�s��=�'���5���^&<
u��w�ҵX�J�(GO��L{�|�����s��x7e�O�$:��&{�Y�F�&���y��j'𶵼ƌ�>�W��<t���n�Z� �o '1��cƆ�z���tq����ϊ�a|��A�8���եK��Ysm)����t=uB5�7���{����إ9x�0Ɂ�����_�9�-^�>z��7>{���V-%y�'��[Q#L��.�W ���m�Jyϼ�s4 �<zf�=	��tG�����&o�R�^��M��o �	#kX.�s"A8S�����s3 4��9,�/f�9<0�[g���[��Q��ь�N���:���@�-��i�r����3m�Y�)n�^F���u���[��G�R]���*���M���~qj��Jc;\�3�=#:�i @W߽�[O^�"�B.����m��y!W���@��&nw�D�Ѷ�"� ��:D�R�Ʀ37�W������w0��WM3��*��=�M�pʠ�c���&Ӷ$V��dt5ze�mX���]7�!�(�
����%N"1#\�!o
?�r����I|YxI�K\������c�w�7��:~���Fj��m�(�[VK����G�F3�%�;��ug���k�[U�mz��o�=՛��:��0�+D�~�D�qU���!�w4:�j��G�t�F�m
�y�����#(@N��@wfH���9Ǿ\3=��4�G�tZ1zM3��&E0���l�oߝYQ�^�7@�+T��?D#�Z�n�h��A��J���mCaI.�H0�VŨ��мP3i�	}j�LbT3�BC�i��a5��Kk(�@D�U�)���M�ȭ za��<�E�z�Ş��i0��z�fF_as�]#1���l�_�).I�^��p��:"�3��bn�~t����]�A�S7�ۮ�P�uַ6�B"�0�y"��(��~@�4\��˝��.Jf����ي��y����d�	��q�Yb��p����0�i�����������i������Yi#eY,@?B1��
9��mY�Y��/��;2���o�O,fj��l?=~cɒ�hQ���I���w��`$�Z�/u+k4���T����7�*h�'/�/x�ҙ���jzQ�:��!��B6MBٵ�M�Դ- mߕ�a�(cN'N9���t3��n�U�:��D�.Q�n�NK�֢�¼^M���Px���H�z��Z: �B1�'۴{��9=���zO��͑�����I�Vq�`�<�L�� 
F܇��l�2�q��A��|������&�/<�;��|�Nb�ǐӛuO��v�Ɛ�6y�,�F��D�$@t�ľ�r^2ū�H�up�����d����매Lӽc��b?�S9��@������6�dF�͒�Ku��%�)��5�42�I�6�f�9��H�LN}!������n���G�o�jV��s��\��W�����]���}a�<)�2��D�>v���j}Yn(�O��2�{2D r:\����p8���
R��_���� :/��F	����,�� MEdGϔ�FB�DM0훦>���jA`Cl�8D�:#2�x������0|Q0��z&&�*M�ǃ�i�;Y`.���.�d���^�3�����>f��ݟ��0X�I��*��1
�`��.���{�Xr�&l�y@-��/K��!^hψ��$�I��]{�3v/_�&�j��<R��7��Ak hԊ	�
������$Rπx�(.	Qq�щ�I�{�$��H���;��! &N�_;*�ބHV��W��z�"�_E�8 � A����^9��U Дጦ��=p�}���:���>̣��mf�:��X�X�I�Á�8b�i��z�3L���@�T���p�b��4��k����F�M����{&��2��Ł��$���n���l_UY�t�眈%O�"��c0���H'�)�����$��FSTm~}'h��]{?(3x낇���r6�G�<̏8Or&� -�Ѭ��l�@J�ӥz�
���W�~C7��Q4��+B`E M�5�1y1���<��<����MX@���#K���{�;Yr��5z�F�NlK��My�݂��8����a���Xb�iY<��dc0�>3��C�Bm�F)^ӗp�Gk�'ϴN-�a<,�������G��Po�<s4������ԯ\kB0���ob\�I�q�]L�P�2!�W���\58x*ڀXeDXV- U�q]�˯'ȑ�� ÿ�!�I1�{4#*O��F����kH�>uZ�wd��ڱ|!k�K�_WJ`��eR݂i�.8�Gw��%rojǎM����
��5������Mϲ�^�Ӏ(�<�/m[.%&R*�g`fG��Ņ�C�>	�Q�J)/S�,[��a2uO�C��� TR��U�`8���C��xP��5��g�����'˪#�a���*1p�-/
��@�r����]�r���$&��Wa�w9��$���q��V�b�:�f�!����!m���>�F��j������Ϝi����td�BM�Wǹ̌(\��{�*��d"�����"m�x��=�"BxjV����g#���7�!���a�uT~E��36��͵K�9Kbh�|G��U�x�Vݺ�-��RE8�[��~9�)����j��yO�m�Y��?H<���G��e��fQ V��<2��Rm���~`V�\��i1��Q_j��>;���	e5ϰ�y�k��u��� a�;E4v�'g"�;w��D�͡ރ��R��pb�Zy�u���7��tR�7�/�ܪĤ#�q4޹a�a,����p�f�2���C�GN�� �	�,L�z���g���Q[
j������p����i�Q&q��f��a�{2�I��P��s�<�b�	zE$,�o�E�J�m�=������� ��-
��xwB���T�I��U$r,l��"�R����e/� �2b��Љ�������e	$H#��3	��&㏳���Z
S�S�`��l]�Mq�����ڊ�'$ž�kH+	��
b�d��Xv�i��-O��/�`ښ4�#�q��uitn]�G��Ȋq�+�m�堇����PbL��V�^=a��/N+�Nߎ��㢢(�fuH�ͦ'Lm���Dߙ�@�vv��v��*>B�_��N���.�+-^pT�-��ܕ��M0�����ViΠXf�G��c�D�v�mAƐ+��Э=`�t�.~�@�!���� %h�G_�I�}x��JLCcJ�)�3f-�0����/� �v�&{�82�#�)���L6�Om؏�rM�����u\e@���>���N>�q���਄���6�,׭�[�����^n�N�Hs�t�޹�|�ʻ��f[1�S�R'?�"Ɩ����+�P�u���y���$�#͙�&���3Ư}#�?�Z-���E�{���`�C'�L� n:�/����0��Tw�h2�JEv�#���󯍄�+�f�f��EJ�	&�9ǰH�Ƭ�s�
�����b@��>�0TN;z��q�L�D�ґ���b�Vt����ji�u��.��b�s%fJ�,�F�Er�G5"���WU d�Vw���58���a�ϥ��*,J��0�&\#Chx�.�q,7��xsin���Ϲ ���QF~����.fU�w��9�ɺ����ˀW��z<��g ��`�y�g���*I3�c�p'�����lh+�f/�rG"���sѰnڠ;K��Y�2�/��or⨏k�@��k3ݏ�<�~_ۉ3���R22ڻ���%4 %<N^�^���ۥ$YQ1=�Ykt�[�j�ܪ��|��}�3�T������{NI��H!��ŏ�"�w'Q�{ �4%V�Mu�w ɫ��F\sv#�kԴC`b�`l�{�Yh��бI�s�d���ݘ��~������
��Iz�Ժ�ٝ�pp����i1� ��B}[�%���&<���Y~5�L����M������?O���������J�Ȇͺ��ɭԄ��TM �s�zmU∛Q���7&���A|��^ ���X��p��\2�m��X�Vh§0m�c:j12��6P�˄)��Z�]��M"�����O�=�a�"j��gP�{��џ���!�G"p�*�ߧd���3Sv�]�}�YK��S�+Ŵ���Z}�g��Ft]>�Q�J� �Q�3�Bu{��7���	��}u�*���
���Ǽ��0��;��k����b��@���ZQ_��������,�d-@o[�Ҕ�h�U:�����_,P�����&��LO)x|A@���+5�H�ͤ%~7sK�m����ڂ~4t�*�Qh���T�|�Go��0-r���V�Pߝ�̘���V�{��ٲtl#Y�.	Sk�P��!���%� 1�#P�4�rL����ɺ����0M���n��L<��?�G�ú��w��b��������#���TLZ�ac>��W,t+��x��o/�]�-�[/f#���Qe���p�@���D��x�^i�\o�&�bo�������dgof����D6�2S�F�E'�v�F6~��W��<=t +���������W/n+E�.`ujؤ�*�+��v�fxC�h �H��G�,ד'�~��!���;��d�q��	�Ur�Q8��`�Ķ uQ�%�����jKd���!59���m"���M$���[���1{��Q6F@�fϞiԆ�W�u����>��X6w_2Z�сu��KW�K1ӆ�n�di���{J��+㊂>;����m ���%��.x�f��5��ٱ㎅ZI�� |�,HFK 秖�3�3U��sW�
9O��13��8��31r��\q�	���4^ D�����`��%�&A�q�v���;�$-�7j��HBKH0`OE���`�h|Ae�����ފ��UpB���9C|l�85gE����;N0݇͔�v@f-��5FEX�Q\�6��yj��lК��e_�|�vC�c���H�jl�21�/m��p���_��/i��?�>��E��+mD�0�t{��	���:��W:�����j��a�g�Ϟv�َ��q��X$���P���nd�f��Eظ�f�Y�ṩC�s�+$����5^N��"�y�MЙ�m�#�`���{8Y����S:#����}~�
p�T�t	r�B澀��!��֭���M��+2�3S	�3��������ʛ���\RA�@�[��}���k��	¯�$MPN^��M	�a&3���HG�}��{�%��w|�._�h��M
dx�?0��}x�]�WFLҭ�rV0��tNuā��gIE�Ȩ���Z���� ���A�W�5�#�3 �+�Z��T��{��[dIm��x����We%���w�/e:��r�(�����$�%��̔�����G�P�}A���0��F�og~�ҙ��9�" j����"�����6�Awҫ�p�L,I��AD+6Ov:��Ų��~c����C[l�h�8��EN��v�N�����L�g'�jX���i�Qy��=ץ�I�W*9I�3]-2�Z|��1z^�бL'XH9��AZ����N�P�����y�����-M'�߫so�����\�QX2����sԕ-%7T�m֑,_����l��@֭'w��Y�[����|0�!��D$Z��a���58�Y�e���G�s�cF-���[u��e��!���$A�8�g_I{����e�_�39�Id8��������Aا�R.
#EB����� "���c���vF
.����}H^&Y�n���Ao�p	�WT14AY���l���z��њ�h���i#r�oF�x8l�br�����ʹ��xj(W"6҇Q��aj}�×x����t_�R��4����G�<�o	T�~������_��P�3��
�:��b3�_1_�f�Ⱥ��[ �����"�a6�cZ�*^�[K��ٌv�%Bgvj�I�b��eW'�x��j�T{E�\{��>�E{c���W�}v/Y�nڮ7	.I�U$vKa�[-���åy�DG{P:��NjZ�n[XS�A��f)�(˴|7�A0�a�3��v7j4L!7�X�I<t.���&Kd_�g���VI�X}�7��IU�ĸ�5���;�_��|�U��/.��X2�ֻj������捝9DV��+�{��#&T��#�C��@����E͛�ui��[Nk�z��a���o��s�<���-Y@��66+�T����7+���x����^��\)���,�Lr����̃�O�]fS�6�>�*gs�wߊO�R/���ػs~@a�0D� ��� ��ލ�n��d� q���|(|A�=b�ؽj8}�G�}�Z<�_�{��7��t��<cK�T\zh�}P�Wp�H�?��J�M��%y�t�p���A�A�Ě��G'w�ׇ8UȷR^�����ٴ��
�\t��d���A��׊���"�s��	�9*�۾2w�j��;��]�7騏|�+?��`ѱ�~Q��C���O<�����7Z��P4��
m��Y.��gf'�|���i@?R�4]T��T�ӏ%�7��{\�?^�Wf2�{焦Zg[]��Czd��;���&ߎ^�fc~��8b���ئ�m�yUH�̫������3k*Ǟ�^r���߹x�J]�E��V(�$�� rU�-����������N
2q\��������|��/�:����&DH�t:�) |�H�\��"�bz}��^N0f�VY��N�n7�5A�� �̊.B��Bfr<�]�$��q���t�)�T�7m$��I7>`�ɑ~�YTG�,�R�b2�!�7���г;� n���%�7���h�>��O�T{�7� 0[�����Gy/]��2�K��@kP�u�7� 4�711���N7_���p��؝�|u�c�w����*<ȇ�t�a�d��x�6An����P?������[���h5���ꬑP����Gl��%��2�B<b���c�����W�^w.=�U�����D  &<<�D��t�<���c/8Y%.���(pi1U�U�z��� ��t_,͋�70v�g4Wi&'�ҡmT�ԢLx�2�:/��%�s�*8U�.�hL���2f�n�Rj�$�gl��a� R=�[���HW�2D{d� OTVL�o���ʭ^���l��(ܠa�z��'���p����-��`zԛ�Z�����*�<����s$�B�BmXK7�̵8zҴ>'���a;��̝ٓL6�Eӽ�W����`+;�_�Q���"�颭�<*M�sj�F`t#G�M���ΐ��59�*ސI�ɝO��<G�+;�3̉+'?�q\����ݥ)�i�ش��Wg͛�KPZh���#T9��ybU�ywЌ��F��\p ��S�,�{� ���8l���U�>�M�m`�1����5�-���A��ϓI�o���4w��i<`i�iK���q���Ja�8�+(btŨ2�,Ѕ��oa�:!����Fپ4^�UndY8zI��F
FG!9��U4� ��z��r��Z��C�˘c����Gw�|O��M��.���f�T�/W���>�$�B<X����_�__���og��zBA�ฅ;��'�������
sN�?�O�Vmc+�DY�D+U:3�CE^@�n�oVAY�`�
�P9�mFX�r����?�'�Xd4�uJ���į�L��+�.fe���uv���1p����S�`��T���;Ϫ��EmTh�Ik�L�'Q�y�>�²�k<a�i���ô�y0}D~'�!����p� �� ���8�p�&ڰ��-���|о�y���{��in?g���_sb�S�U�NZ��;�0$I�.��={]��}�]4��?8�s%n�m�C� ��YP��Q��1d���f�����o<���<�]~�R�W�T\�M(�
���إ'T�_��-�u��E�<� ���.����>b��$t[6X����S��j��~� }�_!@�O���3�K��/d�u`�6_Y;h�.�S0�)'S�*�݅N�W!���6���%����G1�SҖX��Ic\Ĺ{.��w���ٚ鎐g�ZnՑS�qu� M�&���Ag�q�U��C����^5aH��â�h����z��4�#����X�N�����Y�t,��%ts"��r�y9�N]�swM��zc	~$���@���y������)9։�W;�3�|'�ڭku˥�E���u4@��d�6B@�UO��_�E�K�xW�͕�s�E��:���R���:�6��Z��v/,B�	�wrj�=#_R�'�g��v�6}6S�y�J���?ߪ��F�{kn�,1�i��p����?m�B(<�m-�c�3��ݺ�8���b�������0�u�j����� V�Y��I��c�omfi9Q���8h&����C>cмF�-��h��Բ;� kv���x��G��r��������7��}zϋ�ӆ��;E��cC��i$�G�I`��n�pR�8������wNb�~�i ���A�o�����fX���ԕnT�@��e�+V��$�	m|�~3�����l]�.`߯x� ���3��7e���l�݂?�+B
F��{��\f2��eӧ������a��� ���$K�����z�u�r���!��lL�5�9�]�gn߁���E�r��J�n٥��:�xň���W��u_t \��T��P����uR���. J��E�X\��|AG�(W�&����d�bV�Bo��������Y|qo�>R���,=�3dG�jL3Ώ���.(���_4�(���uh����.�> �#�oҩ�%r�]׶Ty�/�K�&5xc��`�������z�0�GϱO!��%Q*R(?��Mk����V_�nW����De��Y�d��i�Ov0wq4� |��&v�X�����<M����4���ȝ}�+>������<�sex�*���P��Ԯ��Z��W�F�P4?m�!�����Rv�0���7���a�$�淫����,�i�j�NG;�&z�5X���k8� \f,�)��>�A���Kv�E3B(��e��-n��=�L�8�q��L�P�x�]����mm��<8�ӗƯ@��z;�U.֯���B�J�ٹ�ɨ稑ϳ���Z F]���|t-�@��W��YgD�5_xr�v�Mi������ΰI��:i��g���'�8���� ]�%'�.�~o��zzXBb�ᣳ�fǙ���ThJ�~!W���g���TMkxجph�'�ZY��Ns��nl��ߘ�e�|31��?�'Q\�l�l�8 /�P�\'��Xyr�[�t^�m�kѐ��F�8�q���0��鷅�����a�|Tw�יC��{r �5�"VOy�P>��kЩ�~h��C�˿����UL [g)�K*��)u�[�7��Qڂ���gB��ω��_wB���Lv�v�6��V�-��"�.�	<�j�p��X��	��u&�C������1��Ks�}��+f�Qj�;�L���>n��r2Hs�Ư��C1���1^�X8�s���lѥ��R-�G�͉�e�I��������#�T�-m�H'<��&5&w��qYJ�d�
T�	o�O���Cqَ�@�T����~z ��v��y�U����`�t>�n�8Ӫ�`�t.�� O!�XV��)�R3����j�	���>z�B�%���9_I�ӕ�u����<0τ�tWʨn�3/�T��Y�2�j�VN�s_�N���Bj�w�C��âf$�A�p�l��i���˟hWx�0x]�RvZtG���9?44L�@���u�Gؗ��)R��)!g��ʹX4�k�n��B�aaK��H����e�3юM�J�}]@�q{b���6�s���5� -֩���m&Z1�+Wqٶh�C�+��t��d/�6�Ͽ�7���v���/H�0�J��� �y�Nƺ��P'஠ok�Jo�2�
���T\��ڡ�C��<�P�c���HD�5
e"�T��ol�qZ\+�#Y�'?�|WI�5�S(��3�~Dw���#?�|�jԭ���k�0? �
C���������
�G�%��}b�C.��4� ���zu��S�~W*��l�iW2�V�ŏ걇HFj"��y�غo�p���mJ	�-����:	6�F��ơ^Lfz��çz�"�D�����z� �pO!����sN�D=�dj��x�m ����\/�X:��봴���"����f�)]e���}�ܬ]p�(rel��M�?��k_@Q�?�z�{��I/0v7Mjl�K��t#�Ӱ6k����7�3�j+���y��I�����X@e�����a}
��%�x�^'�O<��7�V;炷_F�,v~����ۚ���R�W��
�Md �]ؔ��C���ш�dJ����	��z�ǿ��i���!���!3�hX6CG8e�XF�La.� ��ܸiA���NJK���i�p�Py53����R��i3���peo�cW倌S��l�3�� �<hĩ�T�P���#%۩�ܺh�@���K@��[��&d�Y�
Xq���Rt=���wzn]��+�3^��Sb�vme�8���<�`d�tU<�$�US�ph:�J~�3M�D�W��������?�ɮ�O��_�F˽���b�&��WM�:B0��j���N�k�I����޻�۟#E��N��ϓ�������ĵ��[(k.�����b�FH_��V^![��g�r��H�\̽�4���(��T煈%Z�m6��` ����,�U��q� EN����"�G�$�e�����:��[��2��{�1�g��Q롰�����za�@赴�az�+�n�T����3⩈��u����~�[���@�=�g����X�����"�����@�G��M�(�d(����ʨ�cx�@�ъ*���9")�h�+B�(,w~��"�S]����!�ᴘ�ҦQ#8A���0�@y�I�,B���W�k\�a����ð�F�$_�u q,�I`�e6}�3ؙ҃?��3��tR��.���)p�I:j�+����C���鉰���nraf��T��:A���h�a��`$@OH�i����7��@)E��+7�X\�e_�$Rk�Ls���W�y	`�I��s�L����'d;� ��y4a��݂�S�[��2���7�Zj�R�<$j��@4Hb�v����@��Q귮/x,|I�unU�=�=*�v�J�hV�*k�k�cߣ�0|~�*,pD�`2��I=�Tb�N_}��>��2���
��4gG�7m]��F;��p׶p����,k�$��ٟ�`^j�p�l�(A�&5Wç��ESĵzt����S��JF��vI�xD��!�p�&�!�l�4�Bc��FO�$�z�c�N�z1�;�6�ĝI}�ZH͎��P�O�침����N{����b���"��e�#�P�k��,R9^��}��[��&Z���Z���iUL�Py2!W���/5��
���H��C)���s�u�u�L\�,PSm3�����j%���c�F���$�<�c��c���w����dT�3����	���%F�H]k�κmE�~�G���@�@�ٝ�YC �jcM����'cӮ�׷�5�nRƾ���0:z/������C�����^Lg<	o�����Y���ٌ��k7Q�tH�]�fiz�2aG�a��1@��3x� ��_��t\����/���9���]�ʲ�w�d[��������7NQ�ʆ���W5Q����r�eᬏ�)�"��K��j)��B#i���0]|��v��%���u��$Υ)�Y/�~L�⯟��p)��O� q�;1}:/dt�6�]�$��i�G��Z5�}>PW��4!ve~e�d%���ҾK����>���i��Fׂ[Z;h��H� d�]�h������b!7߇��SN�T7p-���LS��E�Q����8��gk���@O,�t�"S��� �-��N�Q��o!8�Ty�.Y�{pU[m@nn�۟|7���G��<��}��}i��{�c~I�>B]������ Mǝ�S~�[el-����6?�Wh�'"�n4 �1�E'&�]�[B������%Q#�Vc8���?�;V��#|6$�����Q�F~�>C��iv>
{3O@�}�H�pV�'���
���=����ï5��d�=�5Ȍ�l,%'�X_2K������j9��xy.�&� �=�iܦ�mpF�5[%��ԆB'��#��1Ͳ� ��CW�Dp�4�6����v.��ܫ}����� ���EUmg��~��e'���FF���� ���R_�xGr�VRU�P;�ly�����������	�j l���{��$5.&��R���H���-��E����pVpg�3�����a "��O�Z�5��kuK5I�_&�o�¼A��QI�{�x���F�O`1�<�%H�AS�	�,�a����i�o����$G�>��0"M e��7���(U]!F �k���qfa��J����L��8�(<��n���X�h_��V6�j���;FZ�f}�8L|�2�G�$~�)yn�^Vx_��T����8���Z3<��v��,��N�P��*�̉�$]�F��V��^"��h�i.���o�u)D�� <2�-�Ί�%��d?o�]���&k%�����/^[�s�����	���(K����S u�*�;���h��a�)�]'ͩ�7-)���9�?Òe[&E�7����%�m��T&�A��ːȧi
�|M�N�Pjŵ*ޯ�eln�P��!6�ﮚ��R�[ɦ�,� ����@ӞH"�-�<{|ʡ�vI
&h��@�CK �h�:���7묣�ӂsD�O
h5eKۤ����4; ��W�G�F5M��0{�p<;#̍"G�{ >b��Q$�ht8B�Q�&$�}͐/
���`����EFe���91�܁��:��c	���v��5F��=j�6uF%�A'|4p,_��\�\�)}~�>Glk��-$�OT��� �juiZ�pС�>%�����#���b��^��V��<�>�+i�)(E�����W��&���"�-t�[L-��7
&��Y�i�d����P�w��o"pV���O���7�X��2���I2�ߟ��͔��:�0C��J�lF���囁�t,�"	�Ӕ�0��?��@����V�&9��?���R�f2k�0S�)�z��[�J�=�Ł�e��Rv��(h=iT��m���_����#��Ս@�.����E���Х`�.����b����u%��� �HΨ#O�{�fd�j �ʪ��v����n��
:5�7�I�r��B���&�AҴ�y��q߸�Z1�`5V�qX�:D	&y�#!"q1��c�}��<�'r��ʽ�̃9�/��w��w��8l"���3��3қW|�{��($k��Y'�F�;y�Ȋ��:�p����I�=�����\[�IV��C�����C@U�#-�KUA��������e�S�����4C)� ��`���w�'�T�q���;��)��������
���_�R��$����L��*GP�|��8³8h��8~	V�F��~�f�����>|c�T�6�㑆`�L��e�dǢ`�t�w���b|�&Zy��F��^eS�!���n� u��\ RT+����拓��� p7�"lr�{L�Ed�T�
��h�M�d����c���^L_����߂a��β0����+��ǲ��w�v 83��V=0�Տߘ��g&���$�^�ȩ��P�*`���EX�܆�R�x$��R�� '�"�'��6�p�u�
�p�9�$�?d�ݍI��	�Ʊ���� ���e�@�\�?�:�5�a|�Q�҉���st��h;ϕ���	�	�/�L�6:�7X�=W�Qo0tO���yM�h�xdi�v�\� ��B�	�ӫ����Q���&j1�fG0�n��+�5��3N��7�1SQ��U��.�7,�.<_W;�������!�y$�����	ӹ�|� �Gyw�x����)%޲�^)Z8A��Z ��Bc�ęh�C�k�kf��(KH����8� ��/I��vH�h]��O�[x�]�ۯ�L������w�/8-���~~����[[G5,�aH��r���YM�R�i%�<���#D\�x\��2�Z���^�@_Ï��m�=Ps]� [�S�aL�����7=���L���⍽m_��W<���UVI���@p�-��Kʨ��׫Aۭ�`�'��c�&���>:���wf�
�v���mk��7W�)׶�~f̡��R3�b��6�w��F�D3n8JDieu�#L&Z���B5,�s�]X ��nNo��\�M�7X
.��E��ӫD�y��u��>�+D�g|S&([��mВ��(��<�`���}l�Q���%a�.�L_J(�ymч�Q�K/k�/��|Z�~����՞]�5�Nq����'��`T�=�[��I��A�s���h3cQ �S�έxf��3��Z�@o����M���0�����
6d��	�]�o����[��_~H�i-�v�?`��ktΞذ��1��Ƒ:���ؓ�O�-��P�`����:�V��\� ]�"(���55}/}@�VK�2}U��|�^�z��$�|�����'����R��� r�-��n%J��N�}o[��9Nh��������′s����������Y�\�9������%Ӑhb�W6m�7�"��s(߿���Z��: =�򀻒���N�j������R]A�}�0��k�~����*�>4���T%��/�,d=��$+^�H8ʏL�;�)NS�p^��kѻ����@���"��H.r��ȘB��`��Eiu�k��_�QݫU�
����Ҳ��p2����5x��Q��e�p����k8ǿ���X���yw�L��A�H+�b�O��W�茂�7Y����� �~�`�U��j�V<C�`
v�2�7�J@�eeu��.e��C���,�.������|�D�[��ܯ��.2�+�C�;ZfD�#�t�G��w)C�J;�E�LT$�a�)bOx���єMj�{C���e]�:sH�F$6�U��Bu60�� k̟�����?R�_up����6��r��R� �<FW��2�<�J��4e*��*�����My��z�ѡ���];�q�ga�����s$Qo�W]��`!�d�h�k�����U����K��I�	��±_�B������+0�U#~���M¬��+��˟��}���W`� �ٌiW�\}����,!��,��:�N�sRJ��)�Q)I��@G�譛�K	��y��\�E�{�qlB���w�h�%�d�#X��Q(YzF�s*ZU����hʼ�q�+V����;�pM�)��zQn/B+�X��=�����G�6���;�hQF�XB��EƬ����d>�D���Q�P� 2ȉ)��m��/��E��k���w�����	c�ݣś�*UT�
h}�'�:��R8G��
�c�Eǜr�4�ŰJ�cp}��v�K���|
TC���:1"���N���	���5�C�2���%߸�F!Le�f�ʩ�$S��r�ml�`c(f���1#<�T9i@8�<�d+�)��˧d���L�9�+g�$��ϑz�5��~�g��l���;Skh�b��l�n��?���?���q9̫�!�ю�\뭍5%9�@�^*nEj��aq:�ܢV`�XC���#�p�����f��X-$w����R@l<�=_wC�Eb�y!��wqo|,�lz%��أŪ��.���*���7J���z�o�N�$���4�s;]�n*}I�?����kT�,��g-S�FO����Y��"f�x�T!s8;V�P���i��
�����xĢ�>���#�
��DQ�8k.�f@����$�[�߯��=��G��=���Xe!�\*X��?\��M#,B����s�ۯ���)�w<����|#���D�rŕ�#į�:�o+|T��wƈ�Fy��#;�b��wRCj��u�k�y��d�$�K(�_I���})��!�|��s�.����F�!�ׅ�ęN�.���J�L����zA��i��iQL�g�˩��q��ܬ��$��2�T,ez�/�?�ڥ�x,E���_1 �ſA�����j��'m�+K��b��+g�p�9�+Yd*��y��<�z�Qo�}r�ۅe������P=Bˈ�
��)�/�;�&��r�A{���Л6�H>�nv(\p!�y��A��s�@�<x�[-�W@��੩*�+�.�d��w����N�E���<֘ۿ�f���� ��̏ A�m�p�5}�wI@Q�e%<5W,��m�b������w?�D��6�Y*)�&���{ޚ�5�$���۽?�;�TovL4��=��3�B9�CQ��H�q�D�*�I��*�I�1�[���7J7���[f-�q�jB��q�0m��V��]��3{9���W"�P.�l%op��S_�k����-lO��ŃN��D?��Dm��b�<�HǬ�R�5Y���l�I��!�6Pb?6�*L�ǔ�����2����h�r��gУZ����|�S�M�xi���RJ�johG
  נ��J���mQ���_	,�K��z�����s�u����o��`{��?̀4��r�8(�^�T��s��B��(�̨oQ]���Zy��6�蝘v0�A�=��yR�8t5�bc��C�HH���j���y��8v�v\|�ȴ>����#z��&�c4U0h����hy�SKnpb�;s��>�"'���0����&.Y*LDʊ��*���1��hՖϬ���̄2u�"�u��$i�+�t����Y�a�!?��_�ZT�3�e}��.y���)��i��˜9RZ ���;�XP%���nR_�V�w"ߧ���Y"G��ZK!��%�* dy�j����Ң�n�)��u�S���FG�6();�RP{����U�t7�8����ڿ�u�k
� ����i����7<�,P9���e��WI��*�s����N\�5�7�7�n{"܊�?Ck��O�V����"*��6���Q���*�� ����)��+I�)�ě�bW���'���1͠/�3�:U�P�J�iuB�s���BY�� y�)&�7�q"x�@��v��>E+���M�xE�͝��m��~�JY� s��5�-q�1`�[�=��ߦ�b&׶�@d���G<�,5�J0������&	�!���D����a<DD#k}^Ԏ4��s�]����C�	��3xlA����J�޾	�:[���Vl
�D�E�F��e�
8�Uj���9�Th�x�7,�IYI�/��V��@�G���CQ�?0����K�����O�Y���[M�A꥽[�3����I���n
N֞�ؗpy��z����$�N�AP�t7i�JC(�ҋG^
_��}BR=@GqX�{�hd������p��о!�vi�~�1�x���+b�S�7�u��G'��K��Jg��͠�=�4)� ���xs��Xm�ᬕA�4R�	������S?��1UY���R����|�N"?�PN��,�|u�j����cv�,�ǣ���B��L��V�%��q#GQ������ �aF�p�w�z%[�R��[~��t����!���~m��/������W��#��FG�XG\	�h�뚚s�]c���S��9�^�?>X�yƙ�E��%p6������F���5Y��(��0��ؐ����uƳ*�Sѵ�JN��E@O�q����1�tX�J.��f���^�\�8��;~�����h�`�y�k�&�y]q&��36�5�W�Ѯ{�%D�e��8J��Qf�阸��)B��>�F��:,{P쨈?�\�ld���1�������cG�x���bNpJEtZ&��-xv���ԩi��-Q�p�^��ƍ"�|}Ts��gk������J>���Yf���ȉ:-7�wx�(�9��@$0�\T�$�u���)���	χ���� G�/��Xk[t��xc|��?�8�e�\�Lqs�r�A\۲Ԍ����Ţ^D���1�I%���#*S��t��:�Ko$z!Su����VHgxT:tǚ�w�+`�2�m���5d�F�>������@rk~@}���['�ӎ��
Z{��:����]w��a[�Ng�l�źH����9��l����Ė��ɛ��_�a'vf y�Bg?�z��)rtu�y/����5R�����y0�M���u�o*�F%,n���O�|�*���p*Ju[�"Π��F��r����n�~bmWl*��s�ߝ��]:s���U����
Ϙhc��B�m�l!�2֞~�7�"��~Y�냈ۈB� 3N��Ȧ��fmk 2æ�������<wpX093O���vX�Cw+��puE��R�W�u�6����]�AD�
k������tjhvŔ9z��Cc o��v#��O�:ô<��qˆ�{Ib#�x˱���!����Fa�`�D���
�/�Dܦ��CP"'ǒ4��%�y��~�K�{�E��,O����aG���MܞN�� �*��CxI��s�vq�$�	�m7��m�ɶ[�����[�����:p�H]�Ə�tT�9�b2��_6�}�����{�����-R;q�bY9�ѩ�&�^ޕ�A�`�o$ׄ��|��!���E�b5k�����_QS���"@����5��
��7�zJT����DK�X�T}��g�k?�th�E���h��JR�̍�-���F�� ��$��	�����Q��5A�C<6���l�L����=�
r&U�t4�	��0Q��⍑͂�@��Vh�O�^i�dN$w���I�x�xE��W�0����*Q��k��,��}v�ŭ��p��)�n1�$˿y]��e�]K�t�\��T�4�3�T�&���/��+�3��>7dѲ��ɌL�k���sT���T�O�������D4�h�h�j%KK�tT���6#�-��5o�jd ��I%���|�.�.��k)`&!Et���"� ��5�S2�����A]�Z�rߑ���G���N����^͂��������+{g���T�K�'/���wb���L���y�����y.��!S�ia�>�(]Sm�v���"��5�!S�}�S&��N�p�]�>� ��	/�I����t�2��D�U&�bWK(
r��}�\]Q	� �y�����{��>��<!`O�o����sr!8-�L]q�$/Ii1��.�^�硱���H�*K�`Ѳ:��JMv�7�J/�_q�|��GU���=�b��Ռ��p^�ң��*�x�-�u�'�gkn�@�ۂJ+?����=l�IH�Z���]�]l^(MgQ�ƨ1��B���H\�S�s'��5{qN��J���*/�!2Ne��`��I�II8f���F�=��r"���T��Ǽ"�}�2j�xVQR����1^�U���I���5/�'N��|qMA�DO�~	]�!�� �8��A����L�_KO�ʍ�$�K�Lv8}�O�I��Fw�B���S��5`��ѝ�DѾ+�&���m�{ӱ/��@4��IO�}��j����W-�VL�p��\��i:n���0�Y���c#��L�?��bՋuzyDl��0���j0�5c�HvA��)҇� 	>_���=�Ct��-���[�F�G	�}r��aᲿ�7D�~�8	P��ƒ:vUc;C�xSRm����"��3[Z�W.Q�b3[!Oo��*�����B:ǆ��ժ�T���l�(j�و�,9�@7�&�:i�/�2DR�(;�%$�O5��BT4R�H��bu�C�V�q?KU��8[��R?��Wug!�M%Z�L~�����zD�Z9�d���wL�����7Du,ю;��z��8�[���6��<�������Q�߃�⍮b��/�A��p"�^���1A����E=L�z��tY)�7(Ě��������1����	��u���K�G�Q_���I��.��`"z��lj�r��Q>�h1���(� m�G:���D߾E���n�l�f �c0�,��amY-��k������z�IN�����L�G���ٻ�;�Ʈ������PV�!l�	��U�?l���kP'�DL�;�A�M���=��?�6�8J'�����^�Uq���1�Y:W�>����6�Q���"6��W�d)^��5�7}�Y������OS|]��j���%�{��--�Q������8eC$�ʵ��6��Z����>�:�n�j��8�8�O��t�W�y��J�yO����vC��r\V���0�x���ikI�w��P��%��ć��XФu�}B(���m���y5�� �T?�P fg�A�Q{+]=�}�����eT�+)w{��K�Fʁ��q]�q�'��� ;���8鉬bE�P�?h�����C/,7�**�#vP}��^ ��;L���G�-:��i����,6��4��W�~1$��<[^K��a΁M�����@}aS�D|�U�X��IbN���|�(�)+��( Q�T͛;�Պ����8�6�z5��)��O��G�E�d��s��`�zt��H+��;�Z�!)��,������[H*/�=,��1][���P�l$�顟���x�q h��Mv���pi�l������s:��}A1�8eu�Bt�7�G)h�g'3����UۇU��_'C��X�{��n�c�ݐG���'�)�{%��1��&cy�M��m;���*� ]?w��䟡�|��9C��!����Z��A������P\�9S#�_������u��Mu�:	�j~X��ibZ|l���4��4��e@�þ�ߔ�KL/�|�bN�h����1��}�/j�ZE����~A���WȂ9IM�ް�v|�n����Ɨ�nL�B' �irΣ��.1�8��;�zps"�p��V �T�7��!�j:f$r��:ts�>e�:9��~F#��W�����}���X�]-M�Px��+'1���T[pNt"�4�`hS�����S����dj��~�;�4Ո��]�&���ig�}��ڊ�{5g)��=���
H�*��6�*��_�W��e��?Ġժ��P ���K���n��a��*�<���gq$������`�/�=4�
a��j>�$p�U$��aHx�2w��I[��*�h?����C	���9�9�	��K�r��+3Bo�M��?ǹ����YHn�fIws�թX��!�&�B���
о�s|��s:�f�����7�t/b+�Z�k�(�s����ɺY}��C̪��q|B��E��n�o���n�h�����P�C��P���>L[*hw��,	=�K3���3����-r�j>��f4�J9r4���Q���B@!���t�z��Q�5������)�A~9�aH>���I�h���6�F�Q@4Ą��SO�
S2���O2��q�=�S�A�2H�#2'�AA����~�}�i4�!8���߽)�>�r�bݲ�27�Pֲj�T�~]8~>cp��gQ���Ƈ{,hI��<#+�7���v�m4HN���a�����N��8}�Jnt�[w)f)�Óvd�M!�Ig�jp@�Ӽ��"���!�DȉGZ���t#uD��PW�Y%=��&����kƬ�'�Q�q�t�G5GW�]�|w{.�h��F�����~x-?$�*�OO����r�o��'9;4;<uW��?�[0�C�����9�9σ���V��<[r��r���BU2Efգְ5\��b�8?���)��J2�χ��π-��؈\\8�><���뇎�$o^d2�=6H{��ࣅJZنx���ԇf�M����՜�3=vsw��luUͷ��5hYX,�ba�C��$�2�r,�)�d�]xD	������E�y0�bԗ�PF�H��m��v�`���c�4G
�b2��K '��i��Q��IFT�X��6�T��D�b?v��h~F�!kE-�b{�/�<H�ɻs��<��D��3�� >�F7g �2�/�������I)c^�}��<t�������Q7��K +c�Ԥ�Ƽ�z��P��
�tҧ�j{Ƣ�+#�92�d�@�r�{��`���
E�6�$�p��I�Ɲj!�ԝ<�GIbv�ci�.��f��w(4��e܈￀�"�B9����{��)l���D9H̰c�f�g�5bue��2�nK�E빂��ϸ��"Qd[Q��x	k�f�S��}��Z�D��	P�SG��TKH�C,4����J�_����-�k��*�L	H7��]� D�G�q��*�����68b��WSIE?��N�=o|����9����>5������6Q.��7w�5�
�|��/I��˻
X��qrݛ��0o{���WڅOpyCD�R�9Rt1���p� ���Ý��S���Mb���<�ț2%�i�� �\����&Wp��51��L���_�|Hګ����I!�+��c�"v�[#$h�`��m �ꯍ����]J.�X��z&��R1���Mʳ�qΨG�$r�o�2tf��w��-۽&���B��������{d �s0�g�� �ʭS��ႇ�
��"P��;��w�fN@q�ѧ����d��KP�"�1i�;����p��#`@d�m]q3eA��~�ָy�N�j&��dϤy'm�Ae��?�q$aG�}���~ڞ�-^Y[H\ݐ���5f´~�wbجo��}�����R�,�S[�u���O��F� g�{~h��#+u�7�.���8?�ꕕ!2��?�f�d/������?��/��o����Ø|mۀ��W�]؅��s�����LfjX���T�)�����H�φ�|�����B
��:��(�a{�d�t��0�!>��E䜐bX�xy��(8�M@8�N1�?dh��B�cu.�Q���A��km�^�p|I�C�8� >�|×�_�;0�َ�14�*DS�8�T�ɧO�jvʻ:��sy��x�x�e�	��d0�
ZOtc+W;҅�$:)v@4t��G+��.5��t)��e�%&��PGO#q8�Cb�u�pj��х���>���P!y��ey�.����.�yy��C�VN�|��mo�����R�=+��v%F�	�BVR��[1�zMn#a6��o�Z}	�)�
`ugH�O#�j��i=	�G(�c∹C�LfO�E�H~<i��bH��4�N�z֙�����@O��v� �
�@a�΋ob�����y�Q��)��7���խ��!a���#^�V�{}&	�ܓ��q�v)vs���g~p���"'�ZcE�#�r���dJMiL�(��B�@�eU���ː^H�q���}�Oɖ��>��p�1��Ѥ�_�����U�DKq]���x��D��?Tc���@98�>�(���ז�l����ד;�Z����g!�UW�EJkW�l�Z���ܫ:Y;Td�� ��>�/ ָ��ʓ�B�� �ePfT��N�*�(���R�'g&lm,<؊������]���J�;�p%j!����]��Ӛd�V1�@T�_��Y�y�� n<]*�@�Ƨ �>���6��s���y��;8�u���@`=Qv���r�����S���@U���m7�o�ôVb�#�Q*��UשCM�0�!%5l@]
�.��ơuc;����ծ��� �(�/�r���n�u�#I-�B]�@s]�_�x.˪9����, N:�y���7�׃2%;��a���6�k�U�V*��$P�O�S�o�xس䎭�/m���s`�ϨC:�A椮V:r�ac�ȫY.s��P���;�h�v�f�g����0]0�e�g��!|�7��-�?=��l�$�޻�h܌�E�J�h4���%u��4m���gmDk�P7���f��'����/��C��2�B�X�j�q��y[:�!e��K���@�p��׭��^��@�LL={G����
���g4����͔�����,��W�ޖ���BTҁA�g,Bj_G;�����MJ��=)2�;L7�\�f��|�6�K!�=����Nln�I���FY<.�_���A���_EF�0�n�֭8�Y��)�@0hy�����E*��H�Ly�s/��ӗӝD�$$V�i{�z�}��Zg�]N,$�e�Ŏ'���v����4 }3 ��Q1���b\'�BM���T b�ҙ+�)�V�|�\b����TⓉg�P�����@�\&�7��4Q�)|L�ܲ��aF��D�9���@Fݠ8cOzT�V5<�'��5V��p��a��~7���Ń2}��Du5�@F���@��Xfo��K���{�QaQ�����2.Ou��m����W$�	:E�2z�Fh/I�Y��J�����F�u6M��I���
"��IB��S��A�G��Xc�p�Z�\�	�IĒ�,E�;wr���m�bK�|sӱŷ���-h�m���{Q1��P����3)��<
���O�7�{ə�_S��h��k#���"�_�09i�ݢQc��2�\9V���F1�V������.�0|bD�� x}:��V)�Z�#A��6�t����vV�0���-���Rװ��������qƩ�+��|��E��u7Աk���#� <wn��V��I7;a����L�������U�i�$�����~��bX�"m���\��
9k�������Qզ&����av��`���LvR{(�����7� ���;g5g�����B^+�V�����f�Յ�����?�z,�{B»:w��w$·�Ц.n�R�ç1Xކt#I�V7�#[��9\�pf�荭��&�bh��$'�~��RYܿr0������ߝz�`󵿔"'��
�`z�}��
r��<=��`i�]�
���nq:�A�$2S�m���f�P@��Պ8B�ahmۡG�n[�(t�T�2��.�VƝiҸ|�1���5͔�v_uF�[2�!��<V���v'�~j2�2q���c��v3�#��U@�yX��H�}��H��|H<��$�3[A�D�In!�� �6S6��·V��m�E+gC�|�6����[�XP��-�o�@w���oP-�2#TE����:�O� ���wI����Xw�� Pe>�ø����	GZΥ\>�Z�V� �������P&Ö� ��2bO��
ɹ�;D9NN�x������(B�I��2�� X����߯I4�hg�I���'�}�I�8Y�*Iy��,L_������d�e_��1gx�E�u�`4//��,>�K��b'��5Zz`Ӆ��x�4�y�X�0��h��;�Æ�ʱ��	�A5[}`D�nT�2f2�X��Td+_  0j��p�����[h��"�P ���n��3���F%ڵ�i�F�� ](��ٳu�q���&���;o����I�]�]���ջӌ-{��:���v�#�L�I���Ψ��%X;C �Ȝֈ�0��^�bp�i��f����k�f[`Pe���Ӳ-�n'�x�7������,�a�Fg	��
����8V/"n�󓼮������7����X�6�ү��6�G�'܃�h5'�����U�W�{�v���<�j\6y�I�{	Xb�VF7$�O+@��>���8�n�s�n-�<��A������Ä�׷���"x���\`�p-�"1?�K�M����%����I��OgKtqQ�^c!�|�N�_5����u˟I�ۥ�T6A�o2R�L�k��,-��L�݆6��m GoG]24,��T��J�[���z:@9r|��]�%N����
��#�6�/��̬��$�!�c���e��t��j$0�8eD�p�}CGl�����,��v3���^r�
Œ�{,{�wʯ4�8�<��:�5��>]6�|�Q>�y�^	��_�i�����S�Hz� *��!vY0s�M�j��ǉ�!���h�-{O�5��; ���P��͇|O��E:�~�eI�"^�=�m�� Of�6��׫[W�3%��φF�i
�-O��1n�8�r�wk(�����P����ZL�U������.��ο\w���V������$��yr���D�u�W?�3l��s0�������;;>�o��z@c�#R��`P�q����l�hn���c���V����>,��n�=�@Sw�����"tqV�c�5"i�#A�X*J4}�����_�P�F����c$�% ������o du`C�g=��۾� ��Y7�MI�.�*���5��)�4 ɚ��nO}�6>���AhJ쫮�;��Tǿ-�CXL��?91y0���ӣj�Y��>wp	��]�^ޜ�J�ú��u,Q�/�:��ok1}T������2/�rD�l���0��d9!�-IWGX���	�LUT)�y���-b�"���#צ���ܝ��%�R���܉�bQ/I���W�Y�wDd�/�
���fQ����9��I��ɜg7b��'�[�y<e�z�/3�K�N>|��: &��#yY������y-o81�N�߻��f���.'�U�/1��YV�Yy�@�=���Jb]��]ru����D#?W�K4�yE�[���{���9W�ΐ�΁={���M��-KC��χ�_5t"��ö��E�F(�4��b�#�,aF�D��$�V��k�A[�Z�3�鷅:nN��� E?��ã��Ϝ���_bѠ�b�w��:��Z�6aVr��ϡ6h�Re��N�A�.��"���r���|���U魎�Q}��B\�E�c-��u�^gS�u��[׊0wLB-^a��v5��}�!}z�X��tV�Ta�k�J���%T��Yv
�,--a�P`��U{���!�l�V�N��W�N`��68��洌7+��8��i�K�J��6d�T*i>������}jr������pI��5��\wT�.ҖB�t,w	Y����Q�z͹����� �mNib����Pܼ��ו�.~	w�l��'Չ���Zm�;Nq����ym�[+4�;h�~���.�!�^�H�vݶ�Y`��+��O��:���@ۭ��MB��.<��~T�{�?fP��S�ZX�*o��^��qA���	��������E��ȏ�m�rY$f�����\<i�ʒ;a�\���SQs������Ǳ�J)���i��G�%�Yrq��G�î���9%����F���eƝ�S�E��$��V�tc�0�їZXZ��w�1~{��%�Vω�z��b4S,:�'��jmÑ��V@ j-�~��AXA�2Vb�"S��#< �">�Kd�����&���X6�ܶ�?���3�`�!�4s2.� �.�l�򝳰D_�ːޑ��B�i?����a��9�a$��$]�=��u�~A�f � ���s:$yr��+��T�U�(���Z�RC����A�i�a}�.���K�Hv�>����b���sc�I���� '�Nϲ�ˑ3$��g{V��.Â��!P\u��+���� h0�\ثy|��sd��!2�C:Z5S�AJ�B�����snZ�I\��p�����+��0�6����>	 T�����.�R�ח��[�>��<��x5f�[k\���e�?󱝅t�8霴��aQ�]�
@�ze)/���
�Qꄼ���iC����&cb�΂���Y_��P|���o��k��nA]�8ꯘ�<��9l�Zh}w<؟1Ń��y@(�Rޘ-��O/������A��w����FӶ�<M�U��K��&�{T���?E\��1��M��L�l%#K����8ܳ#X��U%'��S����Н��1r_�5��m X۸�X!f%`>�&�������:>W$�*׌�a��觙�O�{>�ޛ�J0��2��+����V��o��H����h=���}5�߹h[~��Kd�/lO�rQH�_b��:��w"��*gne�[�p&���e"{{���:I!����*�F*��㰹s��c�5xOm`�Ϯ͉��~P��:SC���D}2�{	 �ae��ɛ�&'1GNjD��������Z6o7A\o���Ԣ���;QS��^ϡ~��9�MǓ�㹯f�83���*�>��>*&l�*�/l���g��O�_�F��J���r�<���Mh�7e�؏�xX��!��� ��!��(��numzRaH~���o��k>l_[Nf�F.�3����1Q�]�qV��5���-��c~�����e�]��#���I�=���0.V��V�Fm�_��צ���*953Gw�EJΑ
�1��w�׷��=u�'8M��p�$0�&/)�����+P��O!�SB�V�=�Y��QsIr룑(�E�gy�"�۔HJP�����Gt��Q01�`��cQ�+����8�} 	J�L>�����Y�k��wdDuo-��ךcGpq��գ�q�jZ 1ȆOSf�Y�j6���:YKaݍ1+���*��?�/�mZ/�Ps�	�W���rK�F�z���`k�j�?6 &9˲��=��c�K�O0x�w/��6o����A�6���g�m�l�plţ�_��R ћ���eemĢ�t1$c�͚,���s�4H��r��*��R�ݓrQ��1u��yXyOM� p˫�MHbh��C�@:�o��B�%��݇�� <տ��Z|�Yn:ɏ�V�`�����t��
By��X1G��}�� ��ֶk{�Jgq�神����t�m�/S�δ+e���8D¶.��+�2�H�T}���+|�����*�39e��d���T�M�楙���7��j,g�ށrw�8#��pF�ͧݘNHu��W>;�b�_c�`07އ z��/�t�m�:� �?�%���Mk��:t�5����9���V��~��q\���f_6�˗I���H���>��9P����}��w#�1�U�u����Qw) &����A+�nQl<=�n����/�wL9���8�@���t`���J�V��#��%t��Y�g
%N5���*0��;�B�DR^Pٵ�؈|�m�	�B(O7�xh���I�3��%��1���Uc �-�<p(�%�eM��b��E��&���t[�M�%Ȼ*����~s���C��f�l�x���	 {7� W��	*�v�ow�>֪)�۠��2$m�od7���J��D��=�R5LztY�X������W�|�v�37��Z���cn���a�	�N��x�#s�G�����?p�A@�^�����>���;��LIO�K��l�"W[���@���˛��NI������θ�w����}��w�o*�8�I�9z�(m��hc��WZ����e�>԰����<��� �ȷ+]Wؗ�o�I���i?0�x�~�ܴW��x���m'A�u-� P�K8���s��FB&F��6X]*_w;��f2荒��N���˿�e���?�:w/��2A� ��q��a��b�����(ܕH"B6�<�Š_����a`�w?i����������D�Ni��3^Y��l+�j��,�,k	^�z )!�aI� ����0\�\�Q�� �X�a~8��c�@V����g&�bE_|I�;`�Q��엘��!q��D=�<3�f�l����Gdu�>�R�!�ȩH��W,���a�Ns�P��-"��r_4�٘q��{l�	޺�U�r�v��nG%�H�1��r���wQkf�|@�^����[^U\;������QuE�[1�ܹ}=�˼4ӂOЩ�pp�r�4��='�L���N�|7x(�Ǒ��z��f��Fg �ɡ��A��vͥjb����
aG_�v��(Z�j�88�E<�L�?܀�{>b��W+���e;�c#WWN���[Rul�Y鐏�`��VR�	��7�'��|h�␹�zP��sL��1C:�%
Y��T��LF#J<��r7�>Z��~$ p��]T=�[�p��\9�H���/~Oc	�(�1��؇�-��q��Ǉ��$�`~���DU��򟐨h�'��Z�`�y�F��L��H��~�ô��UD�ly�rMk���"��Y]l]&%}���!��������dZG��<g�mH��jk��O�Җ��S�����;K]�6yt'�r��|�]egN��KB�$�1V��{�t�[S�lú̲H�f��]���S5���'E�$�N٪�J�;�?L�5�u��
�R�hY:��$.!��=\��t�	#�ym��WD���`��Z���n񏒝����=��3|�_0�f��'�|�I���E��� X��b��b�\{��C;�ug/!�t�P�4	�>�$M���E����kib���c�f�r+��n}�0�D\��ޮ
�Gf�8�P������0�m"S��	�1o�hE�Bj���|#u'eY����b�d|��{�ZXk�fQ���8Hڦ�Eo�w���!Ƿ\f#�{,�Oy�)�T��f!�9�U�i&{]g�H�pN��;;|4�¾sZ���UQTo�=V<�
+��-wfr�N�����y���A{i�M� �I��s"������@[hMW�v+i&f�,tj���5	u5 0+�`����6GH����a��y1:�������z�.t�@�0)+�� �ަ������z u6%q��T&\�ѩn7�B�Q�����a�pͦ���/؂u�^�
P��K����*����9G8����:�Ln=�5�NI��CN�3��w������M�#�[���`��v��8�}<{N{�ȫYm+�.>�.�e���Nd��,�L*<��-_����/6��\�`oj�C�<o��g^��u��Xj ���>�4��G�B1��(u��rR~�Vs����XO�J�)׋�;w��P;fS`ڳ��G8�wV�S�4:�g�9�/��b�%I2���9�Ni?�"�V?�T�]�(��5T^$�9��@h�.�΄I^h�+�JZ���y �A-�KDbw�|�y|�r�⿺��(p��j��'���I�M%��ڬ��\�W��3�Z�� �|4�B�<�S�F/�%������j��
Ĥ�K��5,q��s�˅�iW�6��?Η��ZN]�si� !N��_��]Q�Ü�/��o8�d�tV�~���r3�ѽuؚ�S���"�U?蛄�O>P�;���$5��� j�I���\<����KCjާt��)3>�觿��r�3Z7&k����,�f����7憶qxg%�ߋo�/�)��#�і-T�Ơ7�)���y~>��E$N���%����Ku����]��m�n�f�����Q��-U����>7�@�ȭ�ϳȖx�]��P�1R��z�ꑗ���b��V����3Y4=)�\c�N�J�2����"_����u�xn��=�'��bI���q\˸6�����Z]�D�E�������E;,a:'��~Lw᮲{O���+���TW�JA�O)����5g��(*0jK�&��̕���ǹ{�4��3�	o�V��mqg��(;Z���ې(ݣ���{s�� ���}b�h횞Ř�C�l��O�厂�7B���Z�)�c�����-ym�w2�	C�4�9K�!���e�Ӻ�Au%�<!����,Ł@萔��]��&�jZ����S��Z��mq�$�Y�5�H��k��n��Qh���6�j��B)3�ƈ�M��<,�1�Y�	GI��Pj���������)�����I�p��C^(�wN�!���4;�	�0��"�P�u�`�ț�C��{�+=JH�p���&�
�V�PhxE��v�B�.*8�N�C3�͹0������b�C����`���JjN�&ٞ7�܇���#k7��'���f��N����_�H�Z�<��"6аCXEb��@��%^
A�SFG��*�������\Dd7kܷ9�g��Rt[�S�7F�*��/ź�C�$v�y@�
�b������D}u'r����e��^�(�������n�Y�����cQɩ��`����d�Ƃ���o����Ԭ�{~����yT��(�Β��R�SƁ�~^�)��HLE�姭_gs[��1�j�.C�Ni�'	\�e<q����	!�͚%�n�K�1;f����Y�6��2�p0v�J`.�Q<�eӚ���	����Ǻ+�U��r(�덃i�^�U�c�����RI��Jl�F�MG�
|��Ɂ�&�A���u	XMp��R�_B95��:�1�EfS�2g�!��_�?�#T���#W'�c7�G&{]*�~g���m-��Rt J�"}w8\� �CC=�	m��R4��yL~��Z[��H��bDΏH�d�M�fiE>�WP�>���k�{��B5-Ԟކr(c�_����-.zd)��n�(�ا7�1B� `[�8����!B\�rI�*<�C}�4��� �u6��Y}C�rz�z�h�c�)��*8;��Ync�5�p;{WjMMfe�&�/Ҍ4$���p��׋A�d���oszƌ�<�z�,(:����!�:[SSp($*��Ub� ((����L �3]X�6Djf�%Pt�������B��T85��v*�C�˲8y�����g�����4��"�c�Ym�� L�!�{���5s%�{�a�Q(����D[N
�U���G��Z��(nOp�	4SR��=\V�]7C��io_ѴBr�a�pRH兕w����C�Zh�z�k4�:�Q���hl0L6F�Mw����8����se
�3��h��1[Ci��Y8��Ku�G��L���I���?_���g� �pmcJE��w
�I�1�뷟�(m%�̐��e����&|��1is����#��y����Ge�'^�Υ�,����|5:����G��O쎗hnŬ�8&��<�g�V����19��(逪�V1�<m$�xK �kS�FN�#(@:������Gy	)@dF{0����D-]�rV�}�6�XoN��V�+Q��n�Î�Yg���S�(�����4��}8�c!�6�����ٙ�e.i��4x�l�l@�|F5��Q,������9H;��6%J���U.�����Jg�T�{�������'ltڷ��Z��F���]�>N�=��'"X37�=���*��=@�K�FR��e?ą�`�Y��W�������N��	ރ����9�� 2�D��Ȭ_�>��?�������ꔹ�\j���:���6?.ι"8�0��Zpڎ*��jd#0p"�Ӡ�:�zp����Y)�{łߊ��"�Tp`>	ϯ���[uX�`�h�։
�{ �YfMa����
�Q�g]��)��*�����ꇆi��ٜ�����93�@h�*���R�,F
3�2�d�p[����O�φ�s��J����~���s��A��F\8PE֝�� �t�� ���U�O)�~o@s*�O��
M�uSL��b�������'V��P��w�K`I��8Ą����*��G��}��D��N&f�<nuD�a��sY�\�>�r���A1�����0|�R��|Z�/-V�\T�y��E�F���얋����56�^�tU9�'K�*W�c(���l���_N�"9��,�oQ5���qM�C��Ep��ԡ�I[9U��7��fR�M�S��.�0��Pl�S������U�t�]��s�_�b�>?}�H�U���-�ƫ��:Z�=��@��3��(��ta���zm����b)d0;Ơ~p�&0�2�A�B����W�KT�u�%u�U1>]*Q�0<������Ĉ�v+��BIq���8��ϗ����R0��K�=�i������.s��)GI�]�-�|�(���F�x�.(���˪�,Qq�Ȭ��k����S�ޛ������p~x�M�߃n��T���@J��j�jh��?,���� k	p$n��U�� �T�b08�@�:�,�b��=�,G�˭)Y����È�#ʜ������5ˣ�k��i�gb���չVy�;⸝s&A��h4cb9�G�=�7�툩n��'��t"��8c�i�F3X��K�@7����U�_8��*��&�R��B��z�v�Ⲩգ2��ل<��@7d� z����~c��О�Y4J:5{%����f�_��[��C�t6Ă���[Dw�>�PN��LF!�X�{��ʀ$��5��v~j��t��>����ZrV������?�Lo�M8ڊ�V�̞ީ�����o�0��xu�e�T�	С� �l ���E3���$ǳ��B�4��*��	�"�D�N �c�^�>��C��D'if��;�#R	y���pm��$��>%}>�'����
땣���kkS*g�@�ӚY8��@B��)O krQ]C� ��^�q��3�\g���B̨��A�y���|�5����`؊0@����Nߠpk��H��ϋ���.�S�}a-ytyNm8,;8�TH�( �ݣ��!�a�cK�D{����*��`��8Na����IȂP6���� �&���g�b&�V%��-�����c�d�N�O����v�e���T눐H'�1��L��h�Ѽ�Y���B����'65�X.�2oPS4z��4|�F,r 8>by_�&^XHۀ񏁿�\u��YĻ�2�>��d]8.1����y㪄�[@���{��N$���8�V����ýLP��m�~�1��7x>5�q�����h?w� ���S��`��Rx�oQ-�ܻL�"�M�$cEV%uP<ґ�C���R�jeu������r�h�oְ�>�L�%�GC�k���*r���H |Yєg�K�t9*��2k�3�VЍ3e����knh�<�HB�Y�D�	�l3�il���H��T�������T�+�x�'p�Op�u�g~W+6�)�r<EK�Q-r��mȄ�Xw��.)�)��%X������cD5�T�?�񋗃���E�;挄��@o�������U�sE����G����Š[(��q��.RBҵ�B�����*!���?eH"F��h�x5OҸob�L���ٿ�̂��~���h�����v�Z�Q��bŜ�x&�ɸ^ܦYC�^j׀��ԋ#?:2�tG�e�d�̚$�G� ����/rO�)՜����U�_(~e�0�PZW�n�������j_n"�M�>ZW.6߉�>�7^�a�(a�ͧ���*����� 4D�cOn�����o���ۢ������/H�*h�j�6��3Ƒt����?�Q�	����D�N�O� ���_��]/xV(����b�C��;�<p���t6z�2ī�r+}�tD#b::����3,���W���N����'&����]tɯ_K|��HoR�1�3�;/��kU�#��:��lK�h��Rrro,�ܳ��+��h?2�N����p��E�rʜ����Լa�&, 6��4���4Oa�S�I���H��ֶ�L�ۍ����Eh9�"͗�����O/ɹeֺ޺��?h�ֵL	�o��>�Wtu}�0�O=/���jѫ��;�w(��k[!�%1*�@�UWY��]�4n�u�����\�����Qmat�R'���=���xW��|~�LC��=���&nk����m���
f:Vw�*+$7��@�ƻ��S�[�	�@T~А�s��L'1L���w��w�0�s�|S��D^E��m@ʡ��e�2(�8Q��U�(L���s{Ǟ9�B�f�.'���E�}�YLY��\r5D�0{�����v$�s��$G��PKBo�U���3��w�6�����c�fE!��d������,Jg�f��V��_%�k!4�!����S����V��a��>�B�=�)�9x�I[�v�s������#��&��ӄ��5��ξ4��8�F��K9��/I��߫���24]�5�����b�l���$n�N70��ӳd�M��O�VK�1���1+];XU���t���b���~��»�F�r
�?Ï�)=���L�W�N��ճ���VsD^D�J�j7f6����]#�J�_�kgZ��o
����O��R@����BD��X�y��,s旚d�]�Ŗ��t�f�V���wf�E���?�ib]#N�"�'@ (��V�S�2әK�@�Cs.U��	����'�B7BW٧�ؔ)���Z*���VW�3,�K�&�޲�ԥSNގ]�0�!�Y0hR:�C��L5Aq6�eu��O)�>EO`S�۴��9��U�EA<о�bv�G����t/�)I�N�~j�n�%��1��v��ox���e���D`��)b�V�_؇���\�H�xw�攏���&����'WK���A�����X >ǘ�p�����@�؁�M ��M��>R�!�����]}�:�0��-gGmT�$��쓾� �����C3�^��8��B�}��WG^M^Ճ�T��z?���;��nd���	�Q�8ԁ���J����B�b��<�`�sϕ��È���޳ūC�1�U���x*@��m�K��9Yڛ,|\�	'�C^Խ��[��ʙ���$������f�I����v�M7[��^ e����t����@�&��s�����R�@��.BKQpQ~ŇZ�~���0���@�J��sNq��7a}��_a'�Cy��1�g��kި�,��X�[_k�)���c� SK\�O3�����}�k������8$���A&e"N��(d��c	�ݾ�/�5��e��!��p��N�#�E�"���������	��%E����oM}"Y����;ci:j�p�=��{����@����P�Q�77�,4��~�.H�SKB��\tΠ������s�
 ��]�������:s�R�{�D�XQ���#��Н=tݥ�(�!t� �l�i�����M��W���`�aG4�F���hI�E��kt��9�--�D�������;��{J� �Ә}����V[��2��(�^��QwP��m�S�}�x?�UHB�Ʌ�)��>�����yBX`�x��M��6�/w[�1��|��ƿ&�{e��U*$��3�ZF��+���+�-���]1:<���F���3��ed�.p�)�!l��Ht��K(�yh Bc���|�������b�UP���A����|[:zo��x��L���[��r4\��UFs�̷m��R�m��`4��~���p�~ҫ)���L$����N�AH����H��j #/�U���D�W���r��;=�󡬡�����MQA~������*@{X��6��2�)ZEu_^y���+�=��� ��P����oZO�Fv�d^�S��l��WGN�YXN�z����S�a
M���ƞx�Rn�eẒ�'�R�;^SI:�3yk�@�.Ԡʈ�6�n�w���]3aKo53>�dh�u���cP���C}B�q���ƈ�u�&ۍZ�c�(|%�P1/��O%>X���N�,�a�"J�Ż�(�� w,]��3��M��#';�~3��c�Km��P��>�R?�×��b1�����11�)�����c�����XPOJ4W�{ ���9�`LgZL�\��y/&��O�{�jCZ���9 v�s]��3T%�70T��:̟��v��,�X_|�MFP=�����w�Ԁ ̉GC�H�V]K}��9S���eGw\V���<k8x��+���p��iz��ǥ��C k��D;
�sŕʋ^!��>�|�8Rr���NZޏ�w8����@\P�ɱAѡj3Rә_����c�	����7��:�#�h:H1M�ڛ_P\dT�aTV��"�Qz�ْ�iN_H}�$2.w�r�	UC�o,����{�WZ&�����[N�5	G_}B�y��EDIah׿o�� ����Lq���]A̬��K���W˱"� �	���b*yA�,:�*���o� 	�ӓ
��5�瀞u��#�)���k4��I�L��{U��8,.�=�u�ީb7�9���DFQ��Z}]C�ZR#�! ��	�����KC$�O�b����oO��g�|D�yKt����Ll1V�r���ͮ��]����Nϋ8�Z�N �hzFR\8�N��@�����Kć�?����z�Za��M��r+�U�%�Y	�
��HI��D�q�����d��@9����e3@d���Lc� �Zgp���������Ϟ�q
UB�y�Í0�1�m��TU��p�)���VKZ+h@��Y����.�Zd�x`3�`W2�ud������h˼�As�Z=F�2�9�<GDټq����M֊��k5Ǐ�T>���O���Ԙ3��K�
ŷ���=�����/R*��0|F�\�K�S�I�"�N����st�le�t�k� Z�sB�uо������!������9ֿK�yTqaS����Y2o[�J�FY�H���6+�W�梄<:h⦄z0EoFH��N��l�.n�$/��������Z1PK���!*��H5���%Cy�^M:��i�`jl%�@:�=+�@~����5��z�h�Z���z�X�(
�O�y/L� "4N�*�J2��%�G։oĈ�t��=i~�o���Z�u���d�R��V}���K��}�v:�-�N6��j�9,A��cQ�� '��o�K�o-���?��Ӽl�cD�*��a�s~���K[v�e��OJ#�v�o�XQ����K���/�1�1��I.��s\w}�+��
 ����0�����b�~�x8�U�sq|gsb+��._~�U�͗6W�c�-���V^��YY�V�/ R�U��e�����.^�>��mֿx�qH��/9�g4��?��<M�ŨJp755��tT��$%p�Ye�;�����ً�d]5���D��(�z�����U�N=>�����̺�"ԝ�`���p63�B�S֚:���uo|�W-NHaB�Y\����e�����ش�?��� c���IA6��d�q0g�>�C�uyke�%d}���K��&oP$��%ը�X�O/�p��U]���j�<����i�A�R���bF��Kb �]�:��N��
�<�y��WZ����Ř\��re�v_!Ȯ$G�[1r��6��+�]n�5̤�yb�
��z>��]xGq��:t����{�%U���&]��Η8+[�ϲ��|^�nn��ț��1>\"U����r�M�n_Eo�T]�P��Z}_��)_3�#x\������8.���O�+��(��v6k;�HLjs.��m�]��ŀ�c�Q�Pbl3~�S�nGd�=���Q�kYA���MD�+_�E��Ha�:l�����s\xW�L�qbo�)��~����.�Bɞ���o`*�	Bn��}5��ֿ*�#�4a(��x�s.��M>����i�P�D��?7�,�"̛�_5e�U1�t�r|FY����3��]�XgweR��&�v�P��ؕ<��9�PxMa��	g�2��A���'�(>vk��;�c�Ȫ,��%���9�Ah�1�=��h�!���4T�/ya�͇�3
C��Q��w�K�����wO3���V�$j_���A_�o����n��؟�N�K7�������m'���cQ���rJ��|�W9,؞h�E�����${����Y�.���� ��B��2�Y�
K�єsE����y�(���7I�U��wȡ�j�4zF$���R����΃�4 ��e��؀$� n�ܔ,�3=)�J�̧�_}ɮǮW0�#��h��k�]Y��b��*�2�~IrYΎw\��a�o�i�&t,��
�:��O/�_ӨR�$4�^kÚ��M]��YQ`5�i��%�4��7X�Ԇ[��x�f/6�ݗk�6F ^K�խJ�~^���m��o>���3_���Ѷ�w�P����1ke��m�M����ᄢ1�g��q��͉��h�d��EE(ܸ���`E���` `�6�ҝ8_��b?�Kv/�I8���%�s��n�=)d�W%���?�>ǝ@œ���J8a���D��E��<��72�%�����Ͽ�_��'��?٢dT`R�#�1�QN�2k>.�S������z6�W�ҊpH?��BV�6d���dg3��n���Ҁ�����v�kB��$<�~�J�E�g�$݇%��r��2��#t�$&2�i�H
-?l?�&I6NC.α���E��o�{��e����K
�/sk�N<�������V���,Jp�U�q�Q$�"�N����QpRG�D�Ж�)���OG�M�P�]*��x4�E��0�&���@h�iMJɬ�����0��S��Z_�K���- {�e����mW�GM�i������L=���'|<�����T-�]Zl%�Ŭ��/�G�>ͮ�����,k��k�s��@?����f���۸\�o0�ܗ�'�EZ���S'�I��e^(�|
��b���:ݣ�2ԛ��΃(9z*��%��,�ݗN`C�����=�H��P�D�e��]J ؓǐ}���_�3	B\�N�Jԓ��a�-��=d��rNe*.E��W{��.xÖǆ�{����~���f������t���j��$����pq$������ړŉ�z9��u��V���Zo�5w���h;nu�_A���^41*)�YC`^�i����?ߟ���kc"½���K4�SHD~У=��C)3�4���ڀw�fV[��B�2.�_�~��Ƴ�렐�>9[���B�Ļ����ؾ��P�+zڅ�� `!���������}��[����Cҩ���x�CrpB��i�'c]n���r�h�����L������=4��@���V���`}����	���Ti�ƛ��yG�fr���P>^X�-IR+64��5����EXañOƞ6��R��i�����LΘk�|��`��έ@�����<YH}T�����V4G!�]�6��ŵ��1�,~TcFkb�a�~�06&��\�]2�V1��ة�YQ\������}agʽ�B��-�)mj�4*o����3[��	�?}��{q��c:�?H�'�dk㮅R'��?�<["V��l�ස˫`��v��[D�9kr����M�O��wpE�J����\1��0�a�Q���� <�b5A1_���2��JM��i���Ro�{�=u4�o��[@kh+�X3��4�:�m4<�O�� ��@��f�`���aw1I���{�iR!��t1��>�g|K%���:mx�G��O����r*���I{�S���
#:�~��f�}�}�[-&���e(�m��C[g�&0�C��Y��miΎ�$P���v�[~EvKNV�q�i�(n`4[A Xq8Z���{���m���I��A?U��|ؕ@-�j���"��a,q�&\w���2��e�<S)1��e�h}MZ���@�+/d��8��H�C`�ve��H�
1�nJ���Z2�ޅ�s+:`�_�lԡM3��N�ҧV��(F��<Z��6+��@��X�]���n@����%+o1`�Lք�8�4�k�3��vԑ-Ä�Pq�Wo�+���x�GΦp_F���r�d�4�����O��\)W�IE���Gā����L�%K<Þ_��aM FT�y�76���<�i�^M��-	�P�'��o����Av����s�n��w !m�V���i�F$��D���.(���K���Z+(Z���}ϭ���~	7���� Y�P��?�g�"�R<5�w��CAj�^�T�$������u���� �k���i{�L#�a(�dH���a�u�@�|����~&�_��2���P/$���WKd+ʊ���B=�1'c��m��K�Z�y��9!�Vm���&g�[m�T���c&�Ob)�8c�#��s�G?�����]�d�J;���кT�yKgu�_8n�C6O�m�% ���p`p����=]R��e-u�4�"�Ou����z��TH^2�� n��/SH�����ח��Q��c	��	=�m�n�/(�Rˇ�Jj��� frC�[�9���Jl�4���$h���N�{֮+�#>�to�rX�UD
/(/�Ŀ�c���n�p�qz�F�yYc�f�鍛w���h�ע��y!
)}s�����>�"�SJ���^����J�j-/�L�������ms<I�',�I����o{���[�-n����%���1Jޅ^�?�܆��\@�DO�g������y�X\os�Lryj�J	z@p����Q-7�LLx_���s�=�A�1���ߺ&!g 5-���j���חlF��-�˿�q£_�<�����5H��G�����#0�(y�;,��D�����c��Du�t.�qA^��&sU��H����[T���C���-����S���|2�d7d꯱�3`��2g���W�[�I���٥]�Չ���l�kF�L)����+ԾIZ<@��'�g�/�T��Ƞ|��mG	�
�x$��z&���#���i��Q�<+F*H��� $
�q��Jݾ�\{�̐�`� �� �[���G�)� �\�nt��f=�y��%��Fփ�5�"*��0�G����-p��}]��	W�q�-���R�~��w_��)$q�iܥ:��w$)AG��BRgB˒���yMA���#����H3��2�*x�Z��B��[���KUe�H���~[~�fuu}��`���0�����r\��ז�=]M�
p�P4P��Ŀ%bɉG����Fe���	u��2\Ta��]�uz_7շ�v1Y0t�K����l��2+���'�����@��������=�y�m�p��Ӷ��n��}�H����3��B�S2�ʿ�<�}��M/��.*�g􅯄"W��ƃO",�Bﵐ�J�䰲Q@�K��:�y8�z{Ϲ���X�M�,�Ys�X�c+ծ`<p�z�׽_�"l���%�������r�X>�	�@�EN�f�6���6��qꁫ������4�u8�2�;��vDfx��=fr���ӭ��yz�~���Q�k|��S��<��1����?Q�J&t�������@��ڴN��3#�	�����u��jB����QJ��5������:��t�W�����an���et�6Y���'��?ʩ��XI��fc�V����2�C@����ر��v.y�֍G�gO�
�@�����vy����lz�e�=j{�T����+:�	RI��:�A�����M��*�y`�@�?~�X�so�3\.C�Q��!�+;��x��V�=��8%�т���Zs��d����ԍ���W�.�Ȓ����D:��BȆ�)~`�x6�{Ҝ�9�]�V�J�Pr^�{Ac߹J$����x�1}4�́�����I�5��-n�jw�l��c���\!�"�mIn>�EQ�)u�ܻ,*s�L�NA���mSwXG�L_Ȩnlo�ڛa���q�D���m=�c��� ݄�0d�ݫ�Љ�\�ʲ�-e���#�䤨0�j���?� 2/��H�>���V!������	+2zˑ�'���@F` �2��6����A�7c�`Ys_N�g�k�9������}"��+������b�}Q<Ym�:6�Y������i��{Ýp�%Q�1TُJ��k�n�=8�%�Y(>G36>Z����h�� ��ʾ%��Q*�m^n�5�e�/�ȢP����񀏟 6q1��ddn��o?Ì�Ā�(��i�Ӽ��D��$I8��h���o�R膭��.,� �9箪I�]���]���5�N��P��{��͆��h�'\�|��/F�F����3�u*�6᳟�Eݥd��P�*���q����<�}§��4�A��U|�b�$���3�ːB������^��A��ꎼ%���_$7���K�2;�tk*�r���P6����s�d��ƹ��hf���e�Ss>��|�g��.�ѥ�<����T]���[r@Կ_@��Oz^�^9q�QGE�ja��H�&��GYӝ���Rba?6 ��\ż���5�_Lkf�8�,����@����ձ 7?xqzM�P;\?A�("x����n�w@�3��W�=���ۢQ�n ���W{��XL ��]���>�'�?�/�d^��"5fZy�b�8�M轛��e�������[��I��e��p�x������w��)>#a;0�&?7�Y?����t����'���\�3Gf���0<�~�� �),_��fL�P��zx<\&�Md΃!25)��_�sb�m�5��o�b��IϮ������F����<9� aj�9��}��5cV��;��;���x�e�o�8{�7��%���鼮6a/W=�[�F�C�o��z�d�$���,��N�"������Fr��Ym�I���1ɟ�K6�H����HX7�x��Δ��s�	&㣃�bܠ�9u��*�a:�,I�x����)�I��h���~3�%��t!����,+��h�>��v$�o�!Y����R �"��ж��W�)��c[J�z���Bu�Y�:c� �sdH�*�#ؐ-��fB~z~"����V "U�I(���6�%a�j��� ꎀV������<R�D5ix�u��Rj��x���	�so1_Y� L4���E1V�H���x�t��K��E���\������qٲfx����Cy9�y���ڥFE�tN�r�H,����}�/�Ujzۑ3�bm~��
�l�!��|�3YX��ٜ)�n�(�y�c~���NÑP��m�I�fp">�'�朳�0R�%X��k1tݎ�0(\dl$����fyֈ�=��E���~�O��1�n��4+�����9�BO?&y�@rˬՈ{g�Uؙ�pA��^M�w-��o�Ǝ^a�A��=���&8�Q��D����r���.����C?��!6慜܁x�;�P���{	�=�Т7�6�X:���FW��� C�HD6!?�T�<b���IZ�J���E�-�����p������$�밐ZxVJ�B)�s�̃n��܁���I�v�����
����!;%�l3	��K��mzx��/��p�ta��=D������yL͎�����T/ e�r��1_��L��Y>��p�j�L�՗�-fd��&��zq���l�TI@�[t��!d5`��m:�5��G�Y���$�����������"ð�԰�~]�iMp�j�������b�a(�'�h����}��:��������[��n���{�B��V��u�z��q��^Cd��Bw�Zd�.����w���i��5���?"�J?U6���p|%g��:�����<�y��v�jl������:���}:9����������켩�ݹ����X����/9f�M��P��4QQ?���oO��O��ѦS4����zG��j�$��A�qE��3~�]>�����ù�}�hʴ=��#�o�J��ˈ��_.�]�������gռ�����˶wXd)���O�����h�?>�)m��Sgm��"�:���*LVE�z�f`�E6$�%�:� � [�z@�/W�*J'��O,���B�>��P,g��p�_�5ѢY�<H����`��i� {iMq�B��4��zA�<D<~7�Q%3Vc_����X�A)��Ь�A��^U�h�a�)u�ǻ�|� r��yb{��l�K\��<(D`B���I|��.�՝}�Ӎ���b]8�'P= ��pv�¤�8=C��#�R�gY��Y���0peMb�k���\�)=����M�]T�&�~ۂm�P(�m�e��%�r�L2��by|�L#��߹l���J㎛-rS�y|�L��������̇����+�b|3�v: �C�5�T��6 zE.�<�(�)mr�u_[�#��S�B�h�p�ybP0Bv��JZLZ���{��2��٬<Gb���)�R��1�K>�a=OhR�L�9��&����ReuZ�N���I?�Y��>�R	�j�.	3@bm|Wi6�e���LR�6��	�PwȔ��{Ӏ��Tø�V�!ۘyƢc]D`oY�}�kP��R��a[!�.�E�[d�
��
MG�e�LtXGsc�փ�^>�0�hR&���a��a)��^R"׸|�"@K�m�=g:�BU��2e�򜁃ر7�C�[tH*�wYmY�`�1� 5�������-f����ZU�y�A�I������|e�2Eb/)�/�cJ`�Y�v��,u׏Q�}Akʛ���Zu37$�N�©���v(�e����Fut�����I��eޜ�V5ca��:�� �v��H���?��3�X<]r��nX"��G6�,���0X,)p�\Î7�k���3#��>�&dԑ� _���t�fH*K ׀\3S�@�@*<#�
���Q�&Z��2^��@�o �-�M�SC�p��H~��B�፫l�}��)`��Uu~���� �ҋ���c?^@�;^�ʉ���xBmΏ�j��9�0Áj�:r�Z�K;���1�xԝ�Ы�2�O�Qʚj���`D�B�6J�s�^��v~� |�_���������H���ړ�ԛ���:2Mr�X?H��󉎥�]J
�Α�9��c���w�w%��'O8������� k9�φ~��E�_�c�*���o���_8a5�-y�1�_$�ܒ_�3җ�,��c�X"c\������X1��"̲�1�ʡ���s�L���>��6Z>�?JڞS�u�w>q���O�z�k5��_d���S`{�Lۿa�r��\��+0^��F;p+,�?}�,����'�p���u_�c��ߑ����X�V��6c���5V�,��I���rf@�v׷#�0X��c�Bb� �9ʅa5�i�Żg~�T&p�)r�`��O��Zų�7��"iF�'p��#��+��*�[8`\b�̀�� �;�|b�܉�8����_��ʭ )S?�����-�S�c��i-n�'8X��t-�(�s���<4�W�̭��-EX�w�d:�{N��C�*Ǣ	T���}�-8j+z���'�AF�n�.M�^J�����@O�  �6'�{�� �M��K,�FO?�6��b��-ᓲ�3�i��O�Q�08�rR�h� J�;&�6,? �����
���ϣ��X/�)K-�P�j�Z��t��j��Бќ�8�;w�*mr��hg�%f�OD˚L�1mF�v�'�&t���g�kD�%����L@صSJ��r�cq���>�?��UOp �T%=98���r���%í��p��ǭ~R���<	'�#�z�',0b7�'W��^T��"⧐�����=�(�K��7Wչ��óy�Z��rV�,�Ņ�閐wchE�e�Ң��o݋�&JYT�-�V�]��ʢ�/v���p�����z���"�@�0�P�3=�~պϝ�P��C7�����O/Q髈u�oÔ)� �=�Տ�`e��;pR��Y[���*���0�"FF��6ޠ�m��!=Z��@��GJLX$0ld�0�U\ s���j���+��u��%��0�30�JKZ����7n��\��'����z�xB} �� 7�&��9&�|�'�2��>�W+l�����Y*J�#:ʒSny���4?���� �@c%2]ow�Z���pb���%x�X��,֡�ͣv�ӄ�g�ZHW���1k_~�����+�\>���$��&�Xy��R��Vz����������ZF+�-*�|����I�[�X��\4�����l�lڑ�C�����s�!���EK��� �a�;7%� �"H�?�{\|����� �3u�M��|�ݮ�O'���GN����o��s�h�����t��![[�k/���-	&���=�2��H�Lf4Зݰk��2�$�ʄ~��]�n�1�;q?ւ8�MԾ�����X�����l D�����]�:�?�Y��9.Y:�a58���<��qWB�,�K�>{(#�.:Gn?�M� Jg_X�R���n�Q��!?н13��~���0s�@��`)�
#���2��F%A��~\���V��qS	�����
+^������F]�^ �[��m:���I��rb6`_� �O1O��ޗ�B�~wf��7��2��M#�A��a4�UDk�'o�q������ i :y���ь��/�'�v
�+�BԞ3����_�����x��R�C((�� �h�o�m��e!��m0b@�ݩuCR#(�ΠD�%�����Kdn�(^N$�qB�A�ZM3��);�|H�Q��&�����p>c�Ȯ���eA����O�δ�M[�u�>�)��kH�?:�����,�"�E��ڍ�?�1EmA@����{pP��O�BU�N�n�Y_T)z�s?��?Abˆ�f��.����(/-ƒ�
�/�ߑ�k�>e3I���a����&���3���nlk����x���#X��.�~�8��h���ҵB�l�!Q�U5;a~�O07[F�HA�*M��+����{����_5O�u�����*��#�h#����a₞CO�=2{�V�?#%�'��+ y��Nt�E=+��@�)[���ޟ�����H	����y��_�N�6�%}��u_i5��x����qC����2+�����xk�d���}���pt�No+%ͪ_��l�ؙ�����<��ti 8�P��/	��A�&>��	?]E��yj�T)�KCb(/��Ҋ��c��^E�u��!R5�®�����0���?֙8Ȭp��Fֈ��@Vo؀5����J�Ň�['�[շ�E� _��ײ�� ?����y�8:�?�i�7���1^X7�&իKf���^���w#�ؾ��eRx�c�����[�X6�([fMM=a"QޅH�j��\��d�l�j�(%�	�K��!���	��Y�%ڤ�+�!�&y�����ƿ�����Jf4lp��̈\o[Ƶlo��B�*��Nr��Cx|��e��7���E
��bQ�	�0 z)�Թ\E-�+�AcC���P�~�����������؇��q��S'�~1�������3�a��{K�
��g�Pc�0���+x@f�iBj�VC������x�)�� v
�A�dccq^���PdX�N��S��2�:P��Q��!�W:�i�@	ػN5�v|�w����ZZO�"��Ms����H:ulM�I[Ӫa��'PVVo&���z�߆�l�qCנd+>��l>|�}4}ҟu��0�:������2�Z�Ή�~S�Ut�4���y.��z��\�Y�C�w�b.ӱTf�9�1>T��0�Lj}+#��>q8l�+��4�<�u����)���r���s��Gl���Z�j�`� �5�#%��F2U��?U���#�0%[���[;'{˒%S$�������Kǆ�|>|��[K�CY�MI̒�|GY[� �q�)���4����` ���I���z�j�:��N%�ᐼp����-�=�}-+�vڽ��ᒷ�8�v�vqa�����Q��V?cż<ѻ^��µZ�ǲ~��94�o���'�����V5�"�F"�i�G���#%�������Lw��#X��\�VS��^�^�/��r�҉ݠ�LVMď�RRV(]�ٯD%IEԴsY�=�uܥZg]�}v�3,g-�Mg͙@���N����O|\F٨�T͎���٠t���ꋌ]��˶X�WO�&��7cbB9z��qf*�k�Pٓ.}eIg�|��u��+�@zJ��n&"�=���k�U�ѝ��d��X)�0�Y�t�L]P��F�X��@m�>�𳧬�}���W}z�W�t��x�i��.P،�%� ��3o5mC�Ｔ���Q�q_S�s���Mx#�2\�E�yH����Wm\IʊV�Pm|(��-�<P%&J�X=k.�Yd�X�Q�ñ%#пn�����3��N�Ϡ�����*���:f�����
x��� )W7�>�1�谉#�r%9R�ft{Cg�I�[Ke��{�=_%(#�{Y-���0 y2��M&w���7� G�=<��sI��W�-Ӌ?��)�%���uq��XHd�Qto�c|5S��t�7�������WE&(6���&?�7�?�qTj^U����2��s���w���rW���S�R���[7~;d|�;�#Ej�`\���t��98�m�ۀk�D�3AE��<�~v-��b8��dpܯ�P~��_��i$Wq��1�[�}uA��W�{��x��e���I+�4�BEeUP�D���G*�̵�n��Eh�y+�����ξoo����yh���l���\��BXI�p}9�������	j��U݂�I�E$ե��kC��B�?�t�y7Y�	��c��p�Ov�䯿�P�wC�&uQ��T����*"�ʞ�����>��ݧ�e��T��_�����d��ֳF���%�k��F������/3y���W���1QYW�����Z~r0��edǥ��p�&r��^(;�]sb8`�e�;lW�\	�
�����3�O[P>4�O�W����$�#��U��ю|Ӯ���@��I�<�Ka ;�Y)��f��#����9����pKyݔ~�uOM r��
�_�i4���},k�:�Wnz��E��H��i�N1W�!=D,�wL����sdt'��f'�.�����z�"yvC�w.����I`1d�!�"v�*Z�f9�9;��IXrTcx�^~B��*\��>���5�E�����a��h�D���;
j��Z��'Sˋ��}���RJ� �0����."Y�f�Zf�0[[Ő��l���(Qm�_�%�b������������t��tw7��bЧ���#C6�%r��r;�kܚ�ߋc��ĕ������nؕ¤��
��`�����@l����!�.B1��Z�����!鏊S BkH�-?�2t�]Z��r	��ˎ��"����#���̐X%�C�3���$������FL���C�gs61Y?CpR��
k�m�.�ǃ_ :�����𰛕l?>���]f���-�/��/�G����&�B�*�b���^jI.nB�& �w�p�`x��d�z�n\ʟts����72��~�$mO�}�r��hP��]�Y=��W���~D�Iy�ݢase\ ��5�f]k�ܔ_&Ձ{"~Y��8��>1�哦��+U���eO�����������1JX(!@�͏�J"��UD��QӜ�\��Wq�1-&�O����g��􇉦�4gW$�!Bv� +\w���<L�.�'�qZ�M
�B�gg\�s\��Δ�R�\�z�S����_n��ď����/�j#�j�T���J-�6����9�J���������O��}F[�x���l���v_FX���g����0�`�ì�\{7=*��E���0%���n>�B�$A�n���<��&�?�|�]��&*�A���nP�y�rS��#`�>�˼����4V3�����~c��2��7d.77��y�@��2ώ3�;�K��%��W����m��#�w��j���j{��E%4O9,s1��P@ �r�:��!(I'��*�-xs�C�. "X�c�G���[�u!u�]>[�k����m�l��7��}��r��گ���	%�c�k������o%��[���Q���X�r�ܜVtm�'  �.7nd�cl�&w"O^PGAף� ��.I����R8�EQ��bH� ��	����!���[P���w�O������wu���5�h}-�]�a���A���9��ʊ��7Xr��X��x�n�G�Xw��H[B���m�X,� ��t� l��9:-��K=�>���WhC�'�2��* ���}�K�Ԓ��\�s��$�K��u�ҹ�$5���c4`9�U���	���q�Zv^~b��gX�'[�B��=#VNXr)W�q�~o�x> y�TS�:	���JF|�I�����%H�d���]��������'t��ۯ�)�*?'~��p�7�#���c�,� 9��C����
�IRe��A;�.T�� �iC�a�5�țW�Z�	?t�o肜��G]�	d��)+��cq�/���`�G�_��7
e�
D.���$�(/]�U��%��J�>���3
��ut8yK���q���B'Q��#�o+36�4���T�F�e�"d�z���Ca�+�����J������IӸ�����Ie"j��Z�Y!��Y���$R�Ǯ!���M�$���cZ��a@
G�t6���ぼ��oQb�����nz���&���@,���Ffbg#}2X�g3���7P��\�R��Bw^���{�i����9��pI��hUlҪ��f���9�S�Lr�(����QR���B2w�z��2�c	���i�\.���z5f%���n�um��b"\KE�$W�(P�Ɏ�b&�_����BR���q�qPC��'�n8�Gj[0�֍��|�{ {� � .���8@-�ƈ8���<��㷟����E=(N�"d�l��ڑ�!�^��p��h�'Օi�
Qc[OF,�7]}\@��K�����Gx�t��Y��	sk�c=�vt���򣏄�/�:���'I����J������Ą[�UX���W���/���'V|\��R�B��<�SF�!�z��;���0|d&�Nc�z6>(�g��9��Y���B�J=�$&4�g]?ZdܤƝ�j�j]�b��~:�ǡ��}�V�-�a�鼬�X�%��D:�o{��pg|���r?ꛥ�	?A�:}��{:⋽��	GS�C٣&������V��s������K�����ܦd"P �[ls�$��֍� { ��6j�ށ��q�{D��0ֆ��l����'�O�7⪋�f����#-,���T�[$&9�zLr�1�i��HL@���Yh�Z��� Z��rL�j�D�HEwXk�}�Jc��>�|��S��Y�7z��2�B����Ο?=��Z^}u�|Q���E��~T:����[x���/��F9����6*s�\<IfFڼH  �n�ץ�:*G��zbӴ�v����n9q�����Q��	�<��ؾ���TɐV9��^�gh�ӌ�W��&����#�Pb������,YE���t���iF�>�blIm��b�Z����9u�s.��a#�OJe����'�k�w��'W�qG�翳4�b�[�	2�!��)=�����M��W�q�@�q;�H� 
���Ɖ��è`���:��Y����I�����#y��9��}t�U���=�r9��b�U����	-E#YI�3�"�<7�'��Z�-�K����1��Jhɤ%��Q�8�B�E�f;`��Zl��&�z�GlN"aL���u�kŝ��N�	#A��P��h�j��-�������x��.ϻ��°T�������;���'׎9�R�T<8Պ����`�ț��n4ZƂV��K��f�u��#�0<�ǟD0r2��M5�±AlBΎ=�7��B"K�c����Q*��<Öb	�R�֯�����p��jg!�]�!@MO��3.���ޖ��S��G��i_�CEM����(�w_���_n�f9�@Q��$g�g��W$e���#�z di�*H����V�D(��^�X��f{���}+�1�Rߺ`"��aѰ�_D�G9�Nr�����Q֟)�3�]I��乃	�j�)V����d�0�S�(�c�X�^�g��W���@�Yf��P�sa�<�0�����ֵ�ՙ0 >H����g�C��B��՚�{Ja9��5$��S�{E��%��L�)9\�ǻ4�[�%�#y���%��ҽ)������>S��:^b[�]N��Mٕ��)�F�2٩�G��M4,"�P��}x����+=��f��l��v�D2�s��<l�E�ww�����4��8h~=���i���D�[,��u�����e�Z�q��wO{X��(�șB�*� �v�M�>���S7��[�*�U���D���V�{����ٴ4S[����J?���t�[t�Y&�e���|;9��
^;>��L׺��3���k9̫��`m�Kx��N�ť�e�#pО�p����oǿ��`Tu������+�,%���EwM�|�S�1��(��bX�V�5xi�
<���J�5
�#5�["��ZV�;XZBD3����K�s$��ȹ��ڝ�`Y�ދ�tO�X� Y�$�W���>�H�K\��.����R�G�t9K�X�+���]mE�8XS-�z_��f6�1���|\�
I)�*� 䮦���3��g|�(%��4�l�m��p�n��������	%��g<�� eu?��f��\�C{/�d�Ob$�*O9��r&�,����?2�dD��C� ��o���,���5S��NU��j&� �((^gF˲)z��ȳ2�\�?��R�7h�"R��'�>l-��í;p��VF�+�L�;�v$&�
�+��˄Ó��\�7��sT�k�E;P{�̦UI�;�q�G����Tʃ��ί�H����� ����<�p	�윒l+i�-��a�S�H�Y"WE���P{���Rqk�Nu�zkI������@��7��	��3pV,5^�R;���R�`���2�L�*�_@�mCX�c!V7�Y�TRƶ��g�Xz`�E/���?�VC[b���9 ~�ڙ����z<5������0��ׇ�/��w��Ff����a	ɱ�)ԩ2��,�e���6����ID� Z�B(��#Z����tO��c��0Zr����ъz�������'8�	��2� &���֙��	v1����t��S�I�9G�cRd<�Fn���x�Z	���~	���"D�N�jp��@yWv�?Ȫ���;� 9�$���PƖh�p��d���KSj���ޔ��]��xl��bZ&N6d��l��em��wp:<l�����̀9?إlLBjH²9	s��pƒ��Ӻ���U)|@|���
R�	�^�4Џ!�l�g�J� �ڔ0�^����p�[3�L|8�89A����]t^�݅�|�`��u	������gZ�Ml�h5R�Mcg4 ��5�p�V�Y W�`�p����X���@B\��g����xZ�9=�q���N�r'�C=iO�����!\��n�B?�F����(�-�P7�c&
�|�u���[�׷�SWtt&�m	���+#���'��Y����M��z�S��Of��J�4:b�o�G�F����ۗ��z��&�%#��I���w�5
�@+�^x�ܽE.ô"{���%�P�u�u�4��X �r��A`�)J�a�5�q������cW=;ӕ|-�ާURڅ��p<h���<��Έל���`c�IhbW�b�/����c[���b�V�O�,>҂Nu�GL�ӿZI�@�C�&�(�B5=��m�H�����k,E�'f��|��l���5�f�F���eh�L^ ����䁢!p��ٿ�G?�j(9L/t�������lE���ݦ�R�$����%�g�Z����|���ʷ�Eĝ;�v��բF#+Sכ����e-���Oث8����F��g=��|���F��h$�(4/�|4�K�������#mP���arF+c�e%��{�:'./R�嚨Dxd�u�M���:C�i!/B�}6A'�Y��|�Y���:+��>N�LT)\M��ݶ�F�H�!Ec9�۾��4���C%�����r�C�޳��P1x1o�^����],zb�Y�����ĕ۽SdV�5�JѫM�c��NrlDϟN�������d���92Q��KK���<O׍/���KQ���g��#�%��jN��Rn�6r��ϧ�:���8?�L���(�6noE) �����u�[���>�o�-Bȇ��h���d��;1�-��H
[龰1��fxM67���_����� ��W�OK���o>�*������3�lB����%0�vu�vҕL����I�,cj=:D�]!0��/��o��6���y@'�Ϥ��X�i]��et�n3����o�15�Ɗםu3���/��й<E[g�l�9�N}��\{}�k��d@mm�T>�@�u��n�ᬕ�y�m�~�t��0�}�׵�@�̬q���79ʽZ�� !�]ݸ�n�E�̊�E������s��J�|�t��@�?���|��٦�Dk�T7G&�o��F�eW7oړ"^��/���U86�Z�WE�ى\�I��D�8]��������>��d�A��l�í�j3��x�-��kC!;=L	)$�h���a��}���4
eJBs��ٮXc�\<�[��� �}�dӠ��oB��Q)�íE������3�+=櫠�4�ὰ#��T�af��(�.�j.
�
��O�[�w�p`]����` дl�j�\����J����((�M��Q���.�*��Ÿ����+��E&���N?E����s��B�ݮ�)�䓜�1�C���q�mW%�L�ICy�k�U�)�Y��lM�ړ��_�[Θ�ƹ�����J�0.챈ec��"��mŸ>:���c��B]Hb�����vp�D,�$]��a��م��T�5|��H��J���e�6)D�`r
�֦�,�nR4�E���#��*q��}j̈́�8���T7N ��ǳ�#'��^�M�|��Ь�6<�Y4��y�}��V��!���Š���� �i�7:�_��wG�1[vr��o�%6x�hR�$�2��d�b�۾����;�Ar�Sw��I9a����<�DqO݉�ɱ4�LKH2.�nMdJ-O�{��^�|��&ǿ+�cm�V;:������u��������1��&W��ۓ7�*/�(�%��a����O���:�;�Jiui���{s��/�x�q$���VFl�M.U�R���x��E�*j�����zF��s_	4�9�DU�t�G�/���(��U�M��3 �Glrm)YF����䤤o�򉈞-���p�f��Q/�n
��:t��j��90�\u�8eU��t���ž_�NQ���o���c|��1�m*l�P�Z�m̏�~'���i�U_�VA�Uf�bD1$KP1ʢ�ʏ8��9�n�4\ݡh�W^�������4<&�ѕ�vO,�; �!Y��F����S-X�l�ۃN)ˢ���'���_j�+�7~�	.>�j�J>8n�jo�+��@�o���'�{���������b�=x4�`��;٦�z�F2��է3z���dk
����-��eX$��3�af�n�W{@��A���Pj͏��t(r����"@��MU���S8����ӑߌJ�?��U�Ϙ�0��+�l��j�)��u�B�����t@範+A�w/Jcr1o�.�������M)����V�'m�չc�M�2�:yxel���E��E[ic�'c�J!�2p��nA�-4�>�]nݾ{�AG폮y�-��0X��Lö`�_1��5<��bF�TZm��M�KN7�z[1��cy��NM��Y-=�մ���ܯ�Z$��m^O'����c��fD[;�J�7���>����6W��7԰��yH.�x>�)�E�fV�\+�ޡ���8<W$R�Ɂ{��btRVg?��a��gJZl�_�)�0z)�_C��rA/YTu�ai�Om�6������l&t+�	���$Xl�Pn���f����-�hvm��� �G��bĘ傎��H}���@��;�m�I�%)_�h��Ԯ�ʗ��7CN�L��|C+*�����o��R��i]�\�o>��a�}�A j܄]`�j�JI���ڏ�%Hv~��B��;[ks�b�=g���i_(�
-)�E��@���(ŲK�'!d�-�5%���9�s��A�-�?�68��������cǽD>+S)ܼ���d�X�~6�?C-&f+�$SA6гZ��ji����+�70inQ��b+ݾ7 �z��wj��bD�c���oS
*��{�̎ ��9o��L�ǆ��+.���x�3����Rt5�Z/q�_(�+����<
@�:�R^�{��WJ�!�ߔ>��H�[�������]Zx�[d��������Oh�gءص���D���9?�/�
xr$I⨇�G�:ٟ��L����x��.t��*���D#''�|�� S�c�`�ez�An$���-1#�͑X���~��q�3G=����<��G6R6*�A�y����R%@NPy�imzn�%ĘU�@ՄaA�:wo+{qa��͢g����{~�o<�Y=�	5���tK�Ͼ������C'�9�pr>c=i��g|�Ǆ�2k[���R�l��OJs᩹� �58���/j�-�O�-7d�ό3j���A���,�/��gh9!�����4�y$��7�����򇉴!��_kXh�𗂬�>��E�A��5�vq��Pwv�XP�r��A�,�U�h�}<�[�+B�m��"kp|��tr�������~��?��R��1�@(.���s�tA0�!Y�0�B�-��R](@�ӳ�o��Ca����vQ\7g���5a�Ӈ��w��P6z�Yi�x�h�mh6�V��|�D��͸S��G����V޴$�Vg1����jqØvƸ����]���`�'�?PB�ώ��0�l�Q:��PomI�o�K�F�Ӟ��y+}7ŉ2���I�x!|`����J����=�t(��O��a9f��X��P-Cf|�6�����H�z�)%m�R>�]B�SQ�yOԵU��'�B3���|�L���������G��SD	�p��ɑ�1���,�VN��"�Xm�����n��#�YbǮ���|�]k��(�4� Fg��34c#�@3i8R 4H�(� �����2��O֘i9�w?�?I�O��N=JɌ�����L�h���$������$<HW�Y��8Ov�a}����k�aǦ�aw=~.��+2�_��K�k%�:�������¼ �k�<�k;��WrX�lIiБ�Cw09r�?Q���˨cbk��_�eAr��>g#&9{N9���+{{�'��w�>1k?[ɅV��N�����e:w�'�sd`a���Hq���[��8L��w�c��U�B!�2�&iw.�|{a�T����Jٓ�1gk{�p'�Z?���P|���%!�0U��,�{wW�p,�@�L�[�����Z�����\���8O7�-"ˡoO��E_�IJ�ė��9��l��y+K��'�/J�z�	�������4�o����7E$'r;��<�;Y ��{0,���;�`߻�����jM}��u�|w���d|�&[�1�`��V�#|j��JJ�zx��T��t.�Wv[��a�3�;�^ce��4�|����p���t�����~ڑb/�}Y&�N]��.�7�=6hڿӜ|/32?�ӘJҹ��d�qI%�vq�Tp|LZG=����|x��2FF�	]H�_�VsJ���2	��F)�a�)���GW�������f`ĭE%��u���>�}
�	���MJj(�,�9�������LtINN2�\�ׄ���H@kЫH��a�{<�%^�Qܞ���Ж�-�/�f*	�2�k8u�+�,�#�����R! ���*'� 	��2�-��慤�C�/����|	�H�=b��y�C��D9�e��B]ňm���2-����:��<ե�K���Qƹu���= �����F�+��F�(�z�����5�u���T�j��e��1�O(?�${��y���f}xqfSz��8�r�/A5؄ c�7��/���:��Dv�> �IG���6���XTX�!�ii5���Yh	<���`%R��.�v��%eR�e
*�v���,���6��`dJ���~���|����2��&�^^�Hn���\�VQ���*Z4C���ëB���6��د7��_��򣊋�������\T��}����fٙ�/��z7y��==�aVH5C��{�Z���c�z�<P�\qa��A<%@�*ʋ�������J��#�?b�BiͦMd��s3�����߰ճ��� }"y��EE�	�;ć�3��hBPUU�S�X�/����y�7�}�Nj#"^��$dVF���z� V�AvE����{�D6^a�p�JV��^���ucu�������8���wF�Ŵϻ&��/=(������_Wc��Ζ]��qr���
!��~�#�
?c���T�D˗ٍ�{眭�PP�F���\�j-�Ҡ
T��J��m�~Ն����l~{�hi�v��[i��ǲmY�-#�bC�����j9Z
�o����oV�=-�x�1X�� ��v�]�Ru�*�D��uh��Nͳ���j=�v�w�̹�aM�DS�6���U���O�k�ۧF ������o#	����2N#:���`�/�.��}^.-�%��ꯂ��g���u���|Ez�'�ʤf�Ǩ4ejGPf�L<6۔�w�]��3���7cZ��s^��&������\�����Ln�0�	-������KK'ӵ�^C�˿���K6̈́'6u6�_� �s�6J��`��E�:�C!/ ����c�yd�z]���P��e]U�s�S�F�����j�I&���W��Jv������H+�Eߵ�^��O01�B�c�>A{o������?����04��:!g8����tÞ+���[�7���V>u���8wǽ�Z���g/�4�Oi;�F���'��c��G��
��Õ����r�c�gq����G�q����q2�%��y��Q����z4�N��q�-nm��ÿCI��/�D����V�R����yZpF�Dl��	4�\�pS�]p]����t��ʑǕZ�v4�1>�	l x�TV�A�D���|P͕����z[�8��M�4���m׀�9�I�QS�C��GnJb�>e� 4�
��zj�e��2��,}Nt)�v�Y,#�|,�����1��H��m
q
���<xT�t����	0a�{��������l`����|��6�����nQ��Z2��lV������>չ)���R��͛6Q�����g�C<b��^���K-��c����}�oiIc����i6�H�ԅ�H���;�&bp�ԋ�- � Ch�H(ѓ�,tX i�=:�,�H�Z���
vѕ̋���^�X/���t�\����S$��c�.7��tu�l�g51�	���<���w��y\U&56~����ː���?rBӅ8����/��<X(@_-X�G��Z�By�?����y��)� x������㨰zo�)Me=����݆r�u��X�{�7��I`�[
���ok�W7���^����LaZ}�C�Auw]��}qf���j��<��|� Ǯ#�Js)����jo��?��Hc$��"D��9�4v�IQO� E����޿�In�:1��Rr����i���*�TF��Bb4ll�:�H7�ø<�E�6єG�G������_��=Mw [�䦭�nW�ւ��dmjf���6G�t깵u͔�r%�g��>����}@���o���/��wz}��+*i����^�K"�9�)�o��R�ˢ��Z����J�P瑄6/���5u���������E����I��m�LeC[�#�A��X��~Ǥ<&����t��=wU�_�St�|P}�=�ɖ����5r���7�k�V���%-3��wXg6�'�lN-45zQ�pb�~4�a��05����e�P="x��-v\6A(�7�:���q>�~���4%����׀��D|��mX,��N h�i��o�P��i�^���R;%�l��s����kki�_M�Y��� �'�D��-te�5�]�ah��>�����`{��S���ҷ�{�}Y��l�P�C���I�I9��h�V� *�ސ$C�&��0��3W�E���.�a�l���	Rcx����o�x� ެ�����:�-���
���E ocό����@�n�t���X؝J���|�Iqޠ��xFj�n%�e1�j��|���~�P[���3�M�:<�2Q�#�F����]�t��vЎ�3�{�+��*(ߜ ?���K賹�S�>�mx������>��32
S��v�x��"�����f�ΠF��Ɍ����nO�0pϸ;�1x��Όe���I[{`�E P(!����Lݝ~����д��̼�8�^�k�%�o~ $)�f�}�)��	Dھ�-�G~��4AB�����N&����1&�:�#1˶�n��c�W���1U�Ւ)���J<���R�V�0B����)�L|o�*�&��lo%<og9�#�[Vlt���PC�1�p��1c����>okW�)K�6P������Nt��`�S�Y{�J9 ��j ȳNE���M�'�k)��^_�!892af(��q�sF{�������,s�\%ć[#�X�q!� �+�f5fہ�"���}�'�w;�U�taZ@Yc���hkz�9}������ԝ�7��
��̘O!4�4P�}7W]�/:@�T�2�bF������1��J�ȝ���u�j*��mi?=u����:9I�[���^�|@�����ѧ��ME��(3��r��kws.Y��t'�ܵ�rٝ�Opr-�-��Y1P����%/#/{�������(X<n �$]��P~^���b�4�����{�r ��Y��c�8K�9��y��|�"u�[.@%b�sdI�H�S2��>''�H�S��*���Ȃ�	qe5��jOք�_�,Y��:9;Ƞmi���*1��m��S����W7!��߉={��ReE�lp^U+W��]��~ $�`B|Ä�

Q�
�p���Ni���u��r6IVϘ�Z1�]Z�:VdMqDE��NIgr25��]z�m�䃹ي̛�����8��\J�ġ��P���rmJ��9�Y�J/�2�0*>ˌ(�SU	�� <�ϹE5)�; ��Uxe�l��mNw��i(<�sY��B�f�c�����#��c��zH�-���b�D40O�k��q���z�8D1}&i�<5F5,��s<%H·.sT�0)C���ʿ�gf5�	��m,�c����=`m&�;����+�������S�|�)e4:��+[�uە헝���9��p�L���P�+���]|\0
)����1����u�|������*��.imG����~���!nḁl/��f���|�en@�[���@-�h;PЇ>R.VC�.a$����d�����&�#)}���qVJ��H��!��7"
F^E��c���}��\ш[c�� �Ep�u}�rNU�iI�ق���a�B�t2]V%�e����#)ao?���{��4�"��?z�/�����9˄A�hчd�d@����n�C��;q��i]�K"���L�����#��WR;]#2i�c�"����c�.�&6����ϫ�7�8I�^8q�����+8M�H�@-t�CW��E�<��.1�^�>�Xcr�̓�ʩ.��v��x0Is�H@ 6r^�6���x��l:��� ��o�<�;2%C��t�/%X:��8�Ʃ�JY��e��x:���(�y�9� `/d���mfV�:hwu&���>L̅8U��!�_�l�a�����`d����N��D���� 0�&qM�x�̯W9S*�At�Wc��ȃ��Y��nV�*�p�S��K$k͊X��a��v�O&P��5@+�԰�JNT��"��Ҁ�gŸ�� (��ۍ�m�/�N7��$T�m�=���s ��轂"� ��t���+���R=�u�d��P���>�Ä��H��)]����k�*y��^����F�����:8EtXm�#}�|�k^��z�t={3��ј�T������̼�D[�qSTs5of.��tIͮ��%vO����W1g7�ԙ�P�f���ذ�k��V���&�������S�dqd��w]�����,rզ�Im݅� ��:D�j""�ǂ��niq/�xZ�T�T�w�,l����t�鮃eV���?&ڮr��@71�'��j���|�)ZQZ���*�B3����5��l���0�(5���?�3;�P2މT�#�����g�ڑ��:��7��N�b)�,��p���'H��'FǷB�=/
���>��'+���i�&�>�֜�?�/U賂M���r;ï�c��i�����>��flβ�h���w�?�I0��Ƶ��+�<3	ۃ	h�b��9�S]�����w+�1Ϲ-k$�7�v4K�}p9uD�%��'ۂ���A��K�pTDޑ�O����󓍋	�j�q��>�>��d�T֖2�"��Wk���u��V�ʫ���G~�Za8O��Yɓ0��g�R)X�.#/NTU��FU���.ؚm�m�|��WU��W�=sAm�^�1��3eD�&���s�3u/�JR�Oc��5��2C���Ck���,������O鋷v[���0�$޳�lq�tG��rr������.ZY�vA�/�ba6���7�h���N��RZ.�4����,���L�����*0_�[��Xx���ٯ�BÌ��7� �x���w���>]�[?���A��Lx"�zCB�"M�AT�h�T�ю��K�Ng3�-o�ߗ�^�|_8X�g����\�b�	�y���*?-h��}$��u�1��d����\��̱fi�޿�#�57����.���0߅,��|1n��o���w�e
-jܥ��lu�(�`�Qh��~"�Nt'��^�q���Y?������ش�|7��:�����a�w�
����x)�D�3aF�v����W���|�[1�TP׸��h��kK����3u�/=�ا�5`�R���)�.vʴ,G߆��>��B��I�KY¸�:�{�9 �xg S0�?$���1x���kb_CՁ'��ES[K��[�]S�0�Ғ��b���I��(C�=)�&��a��q|��'|�'��GìѠ��߈�K&��~S��#���la� 9���z��;�8e∖�5�p�	Π,m���b��"�N�p��y	���_3�8�PD>���y_3��3� �B��'���Ud�:J��F��-M���[�����l�ҽG�������y��qſh[��	_�`���@�5\fV�s<�<:�|�`�sp$HF�%�煻q��pr�ɱ���C5#q/䍍7]�On ջ���Iq��u��{�\źr�6x!��:����J��4�`b�c]��~���	i���?�`� �jm:'6��T��}����B!�C3lLHu���킽�a��V���<KvV���Ǉ�>��^)�L �B�L�KaJL�]���'�孛n?9��uu<��A�U��c��٥-R�t��* �.����⦲����K��o���|8�J0��U�~�eÚYl@ER����	I��}��O%��<�H�rВ� �0Ӄ�Z/�v��j+o\���kv��Ϙ��2���	P�u��nA�r�Q�TG�b*2���b֥�K��,?�����S��$.��:E�@�k�?�9A,�������~��i`'� �F?i��!��p�t#��V�X`� 7�s�%
�5b���=|X���	�qՂ�0C/E���1�B@T�����<���r;���zk�Tr|��5�2��bg;��_�z0��Q/�i/l�*"g��OΪ��P��_s���Yu&X�=���6��))S���4��&�ű_�Д�sWA�c�h8�/;t+Ov�
t�m�yG+A~B6�m���!��+��AZ��zN\������,����0!j�������P2�5���S��o���n�B &W�dI�4˧�<"BQ��C����-�;�3e�l� �!�������;�s�f`�E�Q����?Tվ�B�5{G�����m�%��ާ;��c�� ��>
~ʆ9'}�/��)�q�~i��S��;��ݿ�+ė�lAC��O�mĭ0;���'�'�W��TV���H�>�Wq;h��f�c�՞õ(��;�b)蔡1���T���y�f��9x�h؊";n�#��"�ߍ��Pv=�	',o�6N��%%�vճmOWV#��2����A�\��Qp���}p9�.C���cҲ/�H�~�td��֖�{�Y��R�y�Nǔ�tݛ>{�[�<�-��$B�u=�QlT��P6���vf��9�*j�W��Ш�Z��7���珌p�	 	ό�q���8��u��W��s鼶��뉎B� �a�K�ذ�H���FQ�4�����琬�D����%��\���M���g�/ڎ�>�����#�Y���@HV-=�jd�G�����ϭ�p<t�j��[:��z�i�I��h�������^��x_J��ߙ���X(τ�����F�Ķ	�˲�L+Y:�Ӛk��,]����i���j��ac&�ɂ�I���p*��E�û�$�����ޏf����i�j�CH��R����KQB[61�tI?��R)�g��ȩ4x«\{e�]�#^��u�v�y�O�dc�i�j}�cRp��줠�˗=�µj�����x ���v�Zb�ա�I����H����q�6�.���-����d �}��-����hQ�)p�C�d��"�x��@8�A̹-ϱ��Jg�?�I3U9J�-��{��� �oԸ�{Q���@%�jwq��S��3��� Z#,^L;d����z�/�.�V�7�����$�c��o̤I�j*��$>0����p|�w�W��r��w�C}G.9���RZ���l e~B6��\V��xr�pЍ=Ԋ�X�4p�v&t�J�A*�|0MD~/;<�
�BR ���vu`�h�p>��2m��3�(���S�-����哬�r���Q�Q�Dw6�� xh��j���ꅇ��lK���|I�H��r�Mp�`w^��˥~�����zl�4�
�ב@���������X���C`)@����b��l|�ڱ��2�������߭�\�F*������̔�L0Ć���8�_�R���q�5�x���a{���(N��nÊ�F�-�t�^�o�~0�*��h�� �ݲ���R�堵)��#�-���ʯ<ˠ�Wl�P���Jy��� ��r8�*��Ķ�O^��?�/��Zv���6��񡐏�/o�}-�*��T �K��d!<��.�oF%���p���	c��O���𸁥\Ϯ@���*~���NE4,����0U���3չS�e,f�N=��>1��1���Ŀ���9�؟�:�����b�ûH�n)�s�c���bVr�@�����
�^�<�H4��T��i�	���#���4�Ĕ25��z�~�����j;��9+�v�{y�+���в�^
����j�T�e_�rwJ=h�ڝ�����s�^MV;����-��r\W�R�4jQ}x�$��E���R�m�>��F�LP����T�[�m�ʾaA.C}e4o��Z�P<��l��Tz���j�=�z��ה�_Z�H�r �ب�F�?|֪(�54�=0D���*���������1�o����Q���0�ϑ�qe���ol-I�袝H���ZňדDQ�,��G�O3�h���T��"�Z-OQ���)u��������&��q���H����4�S�H3f�硫Q���d:9��d���� Ϻ����^�I����ւ��}9;�� g7�#l}$oo���w��e�"����2t�>����Q�1׿���^pRی�;��|��@9��ܛ'�!*�{���:ʧ>^�&���.��Q��F���#�d�W�~}_��'�̌ Ш��9�o6{.�����o��5
����8�S�w .|!N���t ���:W��F�T�L:��h�v��byk@x����6�5�n�}���~qz߰g��M�?d���7Ʉ'*�Z=+o5ea���>n'L A�����K���
�c�H���A���EG-HR�	�� A�U����߯��z"�����Bo����u��p� #��
�[����4�N�8�G&��^u#W���@=��B(h���+�������d�����^��Q춢z���%���?1��l�Am672;f��:�f�|=� bdc_a�)I܋�������aP%h��C�l��]� �c���9���/���烸�ar_O<.ăܵN�����Ѐ[b/�d۞�
y�Ѓ>� ��ث�V�1e�����{>����%��;+�9Ɇ�{.�z��A�q�ݕ5=� ���m]�!F�(��)j�3�S{���C�ݎ����s�$�����4T�[}����@�Aõ���	�_*Oң�yfZk��%f���W_����j�?x$�ĉZ���jM�lFLƂ�4�?) B
��{�1�鶦�{�W�]Ћїh���m?���A�p�A�p�-���t����P�m�NF�״p�g�,˽���NZ���T���i�w�ɫ:$���N���Z��D=�d9*�sS��i��[��KrHr�z��n����6}2A?&��tím�m�P�=�7�i����ό��	R�ca���ȁAG�`�QQ���`(��\��QG}q�܁�W��{�Rv��"�e��	��-͞�T���[������&��B��X�����Yq�I�Nm-�Iä���B��Mj�dd�O�E��ļ�ƭ&����3���뷏9SQa�?�F�����m1EY!�+�������З^�`֪��b�h���.��;H�c(�
3�mξ�ۄo�W!��������f[���ʑB�?�_�=j��P"ԇɍr��Ӣw|�e��k�	���'���?\;*�E����O�����'���A��:͸I��u>�Q
��$�l�T9hH�В\��%Ze�u����2.���X{�\kp���m�����!ᔿ'4|x�1��� 5�}�^���.U�<����D�~��U�X��{G���8-˷���70=X-���;�B�0��m��Qd��FX��D�Q����¿�c��gE����\�CQY�����W&�� ��C�Ɓ�Ҧ�-(ib������z#�(�B��m����G}���Id���^g�����R9���v8bP�n�`���	1��^��,8��W�#��*�* x-'�1f�~� ��u+5� �'�\����6�8�2J�3���v�$�A�}oR(P��`f���T�9�@��;�长�HXq�J
�/q�E.�iQ]�aM�-��C������WwUhֻ��Z���ȳ�e+�(��,w^ ��G�B$\�J?0����ĞSw�,��b�_G�����G)��9,�A�!楯�1�8��,g�B�>���`���,Y ��=/̑\pB��Sp L�%��-]���7�Xp�vV��Ss���~�h7���dL5�B
J���$�,ο�fL%�k=q�
�W�	���<zk�|��Yx?��ҠS偭�&x#�ʜ�W*��蘻�5��e
������
U�Ó�9�%�c�jj6�,4O���C@�%��߮y�Iܼ��V8{`CFI��=�*�qw������#45}yɸ�=�(۰d����\��LEmjK��[�_�E2����ذ-c`}��T����$����B����3��8�K����F<|8L�%�:cY�V?JM�v\x}EȄ�HP�.��%�c�em�X�����D��Flz�L�������,�~�8aJ�^ΰBg$�L�sж�K��b(�Z$;��+����#F�)j1��S>�/����N�6콑S�~t`M-�����l_LU0G��2�5�,`eN]ɷꃁ�|��Ic���F�h�����E���7�w8-�>!?��ׇʙ�i�G�0��5�7h�ݝ������&Sș��K�P\�6S��3�B��6��7�O:>@�f�B]�ջx��b9=4PQW,�%\��|F��,�E����,�0�I�c��	��QZVN�����|�b!���bQ������o~eA�ϝۓ?TRÕ�"�#_���
��_���*SRBbB;Ev���U�,��.�L��i6�~���U��]��ԫ��������F�심m�E\%��P͍b&����� S:$�"�(����o��.�jO������57g�X��=Q�<�~����u�9]�=5�э&���6//��1�d�}�A��<^qN/�E$�l���q40	��p���P4)mI��Vʟ�56�;D7Q��>��5u4)�nQ1KE�q@�-t�c���,s�G��& ����Y0��P��R��p���G��Gp��A,��	t�3h�'I�?K	��q���`vO���:�1������:�<�ɟ�@o3!�_�F��<����]��d�{��|C��5�աj�i��u�VÚ�E�\��	+��T6޺��];���΁�xB!��N�:x�0����U$��2N+�>L�C���*���]�:��t
�::�;��N�xk�ߟ�Fd��Z�7s�C<M����Eۣ�2�֠���S3�b��_kh�Ӥ�Bٵh���_7n���$��]S�!$4D8������|��[��[�7;e^Ty�hw�������,:W��\����k']��v��p��D�#w�# +	�q��I��_R�G2��E#��ݧQZ,�Tg".���	��/�'�מVS����'@Y��Z��g���թ���82.M���*���!�x�V���v@>>�8�Y&�F��Uc�!���0KV�l��ܺ<(+��~��r!�N�?s�b[,�}$�G�;���;��.��K4��L����A��{�����*�.�Q��c���B5�D�O���p� @##l'm ������#nƤ�o�F����@M���H�IWv�V�w�\���e,z3U,�-�:J�=U!���l
�&Ș�YT�V�D�2b���O�C�%P�1KǷפ:��>HY�$*�#���Y슝��Lem0�i�}σ��J�[������1xQ�Z��e_a8w�]Ca��ހ� b%�K�����z���7����T��{����,'r��kݞL/w�_"��z@j����8�]�&A�V��'��1���@Q�T��|�y��I �Z��Bl�t��g�_����]oN�w��h��I���T�����9AV��}O>�1�G��w�Pj��Ȼ1��^�����|��O�[�u�B��!��e�ke�O�zCTR�8?{�D
�i����I�L6h���I.�xR�����+��{�̨������x�n9�'�
ܛ�����-OW�]�ƾ����kX�U��'�_S����a#"�N3@ �t�X�˲V���G_�#1����6�DwMFեI�=��N�p����k%�������:g���	κ,��¯f��y�%��+���#�x�$�,pŋk�A�k�}�q�Da�P��3'/�lI�8��C�~U�S��!�G�ؖ6��#u�`�{b�{+�����H�Z��_ԒB����
E��3�����y����[\���]!>9$��}�ըF��9�r.�%{�f��o |nH������IêWZ���b�
��bt'B} ��d>���M���a_���{cS���ܧ�H��ծ���7�z��Ţ�rt�"VYqL�:W�t�3$���ݿ��(_�!�$�H�n961�iZ9�g�&$�Ζ-a�5�l�7�]F>��(��j�"(��a�ݮS{�k)���v�Y�O/��0~�<����:.o�A�,�@Ǫ����bQ�Ԭ:x���s��;�g�F�b�?`���R¹S�������yo4$M��JS���˫o��h9��}�2Y�<�/�I<M�����%]�ʜ��q�6�MM�_U뼉����������蚉ͦC�Ǡ?2 ��ޚ�iM���lyq�\��16y����m_K|�Ŕ�Ŗ�)�l$�� �g�Z#MRN.�|�d;�p��ږi\ Q���Q�T����4��c��e��>rA��h�{�o��e�!D�����Z���Q�U�d*9�/�J�N��x�A	���R���ұ�-��]R��{F>.3��ԵQv4X������F޲zgvN0�$���V�ko�uq�����`]?�Y\"-�C�/;l����4'��K"�Hw��!%�<��+=.��Vc YRF�(&9��V��q�*U�y��
�� �FP��j�>Q���h����)���������x~L��?6���hG=��w��*���ת I�)A���_��ǆ�C�V�XG�i��gD�v�B-�o.�Ò���{$�%�\������v)D!�r���_X��.@��0�X���1�i6mD�m58�����㛑�Gkم��1�Sھ�"�l�b�T�����d�.�]�
|�ȇa�6|��p�խi��d���{�Ƈu�*�K�!t���u&`��/�Wk�7��.���G�Q��$�j�ݷ��Z~z�Ϧ�N:<XI�Qn>�JM)�Ӷ%� ecqD)�Z�P���Z���c�H���=�b��9;� AD+�0�X�YaQ�g�m�Ь��Z���$���g-7z�<�ֳ��V�������.�C	΃�7�a3@J&�#T�r����z= _����p��L�̄�]� ʶ{�(�Z;�E8����׼n�L!|5X i�Rk���7z���C��b)kż�+C	T<�h��.δ9ݛ��D�����)�셜�ԡ���XXf�
���U�	J3���q��%>kq�K�@�.
�囹�n�M�]x��&��n'K��N S)����F#�t2[�I�]�@i�Uf��j�O�+��g�>����ׂ��YD
��j���ۻ��Li�y���Ax%e���nnF���^�4���,d	����eLL����kkžBك���;�%��la�ݤ��Fz�z���u����*�^�t�Gu�ܤ�#�����ܶw�n,��W!uL�ꂂ�!�{�w�gdr��P�I���\�h*^q����м���'�X�?%qu��F*�d��r/�`����c��QFex���-���P���2W#e��#=��7c�jB��[��]��I J�Lz�N�%�MY5GE����:y,m$���V�2����i���a��@�ҙ���X���b*��`P`V�Dk^�H�d�y�k��H1ɒ���Y�>��Ј������җ�����k��
�Pb�V�6�/��^��"��@���9K�H󠃄���܉X����XoYE"gU3��'O0��?;B`}���Q��#B"Phi�w��M]%F�����������;y5�[-�2��:����k�ԭV���14MO^��8ͳ�r�u��q(��{�#K![ZPGn�!v����$��
S+�"L��d�b4?� ��ځ4l�r��V�yJ���HΩ%��?��뎡@�� ������۟yt����� B���.�U
f�ĉ����6L��͇��L��a���-��Y��nY_�D?}Ψ�ƒV(d�Kt���'���e]�ʁ�-�0�4k
+��o�@�1��BƑ���$3 ����?��@���[�G���S��ʏ��D�V���{��.�!L��l�އ̊V0I�Pr��>��mw�;\�`c�N`��x:�@�@@*�_l��?�5�KZ���!n᫾���z�/�9?���s�Қ��Q���������E�Y����X��(�vK ���*�4�1���yp�,Z�QS㦲˯UK�7�ܘ:S!�x^(o���um���ّ�T�Z��ن��\U?�M��y���LUTu���Bt�؃�5�5g	U�g��̋H�A{
Hɇh�\q]�R�L�/���	5�d>:߸+�{��_f,z�_J�>h��hc�F��0����=F����O5o���y�qK���\�ID���&��}a5���G#��b+�ª�W9y��-���{���yw]a��Y�7`p��H2���`��<�a+K����\#�u$���^A�"W�&2
E��t���	UB�9�!���nY�x�爊�`��6�Q %���o$u��� ˘v����k��~�f�0ּ��޳�g�*9���$�|��'��|K�Lr}sJ��<�n���{�f�Œ!�,�FA9�U�y�z#�r�
�`/����v��wẍe�0~h�GO�V����~ 5�����A��M�N���j�^���ѝ��n�~�(��4���:�Nj���Z�G�������{���u���>s��G�`�kٖ(5
F�Z��N�mF+�7���W��0d��2eu �F���p�m�N�r�oO���������b����&�-gߦ�G>��5r1���l��$��A�`����̹��׀���KNk��H��}�V�/���hv�c\�b�:1LX6���e{.�ܽ�G�X��č5M�*���]���t���*y�%wO�Ῠ6�7#ka��p�m�J�6GwG� ���H�\��l�&����s]�NmP����nd���4K�|m�V�
)�Y�py~���3[`z^��x�'D{��t$�� �lucm�R� �Mӄ6������;�[��8�	����:��xNus�����$+���� ;���Ey=R[�[�Kv��N��.����f���3��wm���F�(�T>����nOꘜ.�x䈊������i8<1L�"z(1����K��Ѣu�Q��i��z�r�&W��+V�@�R�t��`�~�Di��}��Y��j�D��hѹZ�kOU�+&����e�	qt!���N.�V防w�x����)�)*�(�Pn{+k��8��mcЈG+���t��/��g�����ye�gA:�lU(�-c<w�2lD-f}'�%.����K�n�X\�w�VH$1��p�7_��>$y]x�{k��D�V+`O�UVR�\rd;ooL|��gPorGa2�4]���:Z�k�ۉc�\Ng��aD|���k��xY]�v�G�@��_h�{���'�Ƽ`��#.\|��@�9�<4�8�ģ���e��A6�Zd����~��7�����P/��X�R��8/Zj�YBA�ZJ��ܺ�G��]�qIR��\��Ԕ,�(�!��
�]�`�Xp����G��AA_Gs\u(�����a��w��e�O�$�[3;�����s[�֣��ո�Z@�LO��]C�v��9gV�M&�Wh 	�_��Lhw��m����*TW̔��O���^KO;J���	-�tiD�K��d��^
����|�0��~Nd
��7��`w�X �^��C"J�mJd�b��b��������[W-� E#w���mcݕ��~�*w��ݧV6*��Z��jP|"���4�J�`������K��<��d���P]	w{Ug�RE��vv;8�J�<���da����i��Z�H�>���D����:������V$���S���7����S�A%h�0e��U���;���@��_��f�I,��#���}!v;V�G�c����p���`����'4�I�>��>�=�M�L�W�D7g#���h�·����Rf��U;����ܐc:`r���}��D�omz\���[cÌ{=rb�$��/!D��&~�;�R�T�m�Up7��H�\X�p����[��}��"�L ��Tй���v���5����qDg��c<ԸO4���Z*F�[�a�68�V��n�XT�Hh�Ft�L�Q�D��Ǯ)?R�b�}r�)�.DR4�d��������"z����{G[C������>P
��������X��}?�s]�ѥ��l �w�_%�<n"��s�ں<��c���~Y��}yW{)�4�5d:K��E�Ԫ��p���zB��*�;G����,4���џ���k��sH�A����>� /q�͔I��Kx��%��rr��{��׸��P�Ԧ���O6l�x}1+D�|����F�� 9V C����X��6�hJ��X�!���L�6�;=:����w��G�8Zx=�&��ZF�O7��b*# �N��Z<�V�fJ�Qv�e"����`/�Bgjg@�"z��6�}�*���y�pPK�zv��~���(x_�{QHp�,o7�ߜw�\�)����/§fm���0
����e*��=��<h��-��m.����t{�������s����׻,�*Ɉ ��f�ڙ �	�5������$�z��G�?k0<E���{\��sYg�E1�� �fNͤ>T�5��D�����'�2`��(��R-�͞�@��x�R�Y��Q|%>"6(��~Y.N����� n$ ����+W{�9���I��)����e 0��ݲ�@��Ǳ���4�t<B�I!g_Z�_-)�?�~���Ҧ�a���ll��1�՘5`��L0��9^�|6��:�&Y��*J��~H���q&���sC.�%s�"7�P�|��8�ýF�i�R�V���Z]«ϼ�[���T��U%>��i����Q��C��P��_��Q%."���c�٘򄯌���?������J��q�HY�7�.�%�J�k/���6���$���� x�L*Gm�: }�k'���5��Qզ�]�~�B<x�E���s�h<D7�]��Ӽ�l�A�h�M���v�ȍ�*dA�����{���"�������X,3���,��)G�'&���!5�����\�]��}�ϫUF��7��\�!�r�1��E�2ܶ4�$q���~
��������(�ò�S�;?���lKrH������S��8�V5��w�����-���
�V3�}Bf�%,�`RX��dV0�w��4�{z��	���x񑎳�M�� �=��sش
F��F�ۏ�U�g�q8S��6GN�o W�x���c���H��5�|�2�
��t�O�����r�Z�Q�P��n�t��	�~�+1UH:$�	���	��J�:ZFgD�.MU�m����Z��IEՁ_z��aVSsך҇[o�R���_,s�#�YC-�v��^Sd��]p��� d�b>��k�����qh��Z�Ew���� ���<��<�`V��љ�o���b�n�x�)8bB?�(H��_�(KT(�$H�������'�8�;�Hi�_���6��<���l�Sm�T��,�T35�_H�����{����s��46܌A�B��1�i^zb�QOĐ$Q\&�5@�,�j��
8G���]Q�Ubv�.���v�?
�o#�w�]�M�i�j�a�Xa�B/�tH��۩ߐ������w����+ �l	���2��0#���E�F���q�<��v�X~��ƨ��DV� �L������a0���t{+T�h�$�SV�AE��[eX�>f���q$Q��"�qt�)�,A��E��1'j�s� x$n���A9Ġp����`�~� �g�ق�Jx������\[�,}Xs}��QIK.P�اoE�R|��[���#�E�\:zM�.ѧ���/D�:�Ъ���	%�+U�'�;����W���ۏ�M�/,~����/#O� 3kٌ����TNo)s$t��Ur��vO�1/�lz���yE^�2K A0�6!��f�p�G���q��uޟ��'C�]�'8F�e̷�O ŰS�1�s�$��ۊC�tl೨w۟����v��Wꐈ�ZQ�z���~���c�E��eq�o�;�H������
�>��ۦZ�{)�^o΍�(~ݻ���mV>1�rA!��:�R7VVe�$�'���ȡ����,��2���O��� �w&�TE8��V����\i�K�D�TU��|`�8�!w�J�Fl1����	;�tN��