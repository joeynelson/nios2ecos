# ====================================================================
#
#      nios2_tse_eth_drivers.cdl
#
#      Ethernet drivers - support for NIOS2 TSE Ethernet MAC
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2004 Andrew Lunn
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas
# Contributors:   gthomas, jskov
# Date:           2000-11-22
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_NIOS2_TSE {
    display       "NIOS2 TSE compatible ethernet driver"
    description   "Ethernet driver for Altera  Nios-II TSE compatible controllers."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS

    implements    CYGHWR_NET_DRIVERS
    implements    CYGHWR_NET_DRIVER_ETH0

#    active_if     CYGINT_DEVS_ETH_NIOS2_TSE_REQUIRED

    include_dir   cyg/io
    define_proc {
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_NIOS2_TSE_INL <cyg/io/altera_avalon_tse.inl>"
    }
    compile       -library=libextras.a if_tse.c

    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
    }

    cdl_option CYGSEM_DEVS_ETH_NIOS2_TSE_WRITE_EEPROM {
	display "SIOCSIFHWADDR records ESA (MAC address) in EEPROM"
	default_value 0
	description   "
	    The ioctl() socket call with operand SIOCSIFHWADDR sets the
	    interface hardware address - the MAC address or Ethernet Station
	    Address (ESA).  This option causes the new MAC address to be written
	    into the EEPROM associated with the interface, so that the new
	    MAC address is permanently recorded.  Doing this should be a
	    carefully chosen decision, hence this option."
    }

    cdl_option CYGNUM_DEVS_ETH_NIOS2_TSE_INT_PRIO {
        display "Interrupt priority when registering interrupt handler"
        flavor  data
        default_value 3
        description "
            When registering the interrupt handler this specifies the 
            priority of the interrupt. Some hardware platforms require
            values other than the default given here. Such platforms
            can then override this value in the hardware specific package. "
    }

	cdl_option CYGDAT_TSE_GET_ESA {
        display "The name of a function that sets the ESA (MAC address)"
        flavor  data
        default_value {"get_mac_address"}
        description "
           The name of a function that sets the ESA (MAC address). 
           Signature is void CYGDAT_TSE_GET_ESA(unsigned char   enaddr[],
                               unsigned short* base,
                               int             irq); "
    }
	

    cdl_interface CYGINT_DEVS_ETH_NIOS2_TSE_STATIC_ESA {
	display "ESA is statically configured"
	description "
	    If this is nonzero, then the ESA (MAC address) is statically
            configured in the platform-specific package which instantiates
	    this driver with all its details.

	    Note that use of this option is deprecated in favor of a
	    CYGSEM_DEVS_ETH_..._SET_ESA option in the platform specific
	    driver."
    }

    cdl_component CYGPKG_DEVS_ETH_NIOS2_TSE_OPTIONS {
        display "NIOS-II ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_NIOS2_TSE_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Nios-II TSE ethernet driver package.
                These flags are used in addition
                to the set of global flags."
        }
        
        cdl_option CYGPKG_DEVS_ETH_NIOS2_TSE_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the Nios-II TSE ethernet driver package. 
                These flags are removed from the set of global flags if present."
        }
        
    }
    
    cdl_option CYGDAT_TSE_MAC_DEFAULT {
        display       "MAC address used if none in flash"
        flavor        data
        default_value {"{0x00, 0x23, 0x23, 0xaa, 0xbb, 0xcc}"}
        description   "
            A static ethernet station address. 
            Used if this is not an Altera Development Board, or fi there is no MAC address found in the flash by the MAC address function.
            Caution: Booting two systems with the same MAC on the same
            network, will cause severe conflicts."
    }
}
