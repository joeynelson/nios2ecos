# ====================================================================
#
#      opencores_ethermac_eth_drivers.cdl
#
#      Ethernet drivers - support for Opencores ethermac controllers
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2004 Andrew Lunn
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Gaisler Research, (Konrad Eisele<eiselekd@web.de>)
# Contributors:   
# Date:           2005-01-22
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_OPENCORES_ETHERMAC {
    display       "Opencores ethermac driver"
    description   "Ethernet driver for Opencores ethermac driver."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_OPENCORES_ETHERMAC_REQUIRED

    include_dir   .
    include_files ; # none _exported_ whatsoever
    compile       if_oeth.c

    include_files include/oeth_info.h
    
    define_proc {
        puts $::cdl_header "#include <pkgconf/system.h>";
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_OPENCORES_ETHERMAC_CFG";
    }

    cdl_option CYGNUM_DEVS_ETH_OPENCORES_ETHERMAC_DEV_COUNT {
	display "Number of supported interfaces."
	calculated    { CYGINT_DEVS_ETH_OPENCORES_ETHERMAC_REQUIRED }
        flavor        data
	description   "
	    This option selects the number of ethernet interfaces to
            be supported by the driver."
    }

    cdl_interface CYGINT_DEVS_ETH_OPENCORES_ETHERMAC_STATIC_ESA {
	display "ESA is statically configured"
	description "
	    If this is nonzero, then the ESA (MAC address) is statically
            configured in the platform-specific package which instantiates
	    this driver with all its details.

	    Note that use of this option is deprecated in favor of a
	    CYGSEM_DEVS_ETH_..._SET_ESA option in the platform specific
	    driver."
    }

    cdl_option CYGINT_DEVS_ETH_OPENCORES_ETHERMAC_TxNUM {
        display       "Number of output buffers"
        flavor        data
        legal_values  1 to 126
        default_value 4
        description   "
            This option specifies the number of output buffer packets
            to be used for the opencores ethernet device. A maximum of 128 for
            receive and send."
    }

    cdl_option CYGINT_DEVS_ETH_OPENCORES_ETHERMAC_RxNUM {
        display       "Number of input buffers"
        flavor        data
        legal_values  2 to 126
        default_value 4
        description   "
            This option specifies the number of input buffer packets
            to be used for the opencores ethernet device. A maximum of 128 for
            receive and send."
    }

    cdl_component CYGPKG_DEVS_ETH_OPENCORES_ETHERMAC_OPTIONS {
        display "Opencores ethermac driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_OPENCORES_ETHERMAC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the opencores ethermac driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }

    cdl_component CYGPKG_DEVS_ETH_OPENCORES_ETHERMAC_FLUSH {
	display       "Cache flushing"
	flavor        bool
	default_value 1
        description   "Flush cache before copying packets from/to the
        ethermac dma transfer buffers. If you have cache snooping enabled
        you can disable this option."
        
    }
    
    cdl_component CYGPKG_DEVS_ETH_OPENCORES_ETHERMAC_ETH100 {
	display       "Initialize MII to 100mbit"
	flavor        bool
	default_value 0
        description   "Issue a MII sequence that enables a 100mbit link "
        
    }

}
